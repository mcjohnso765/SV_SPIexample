//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN210F (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.


//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN210 (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.


//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module AN211 (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;

           and #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN220F (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.


//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN220 (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.


//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module AN221 (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;

           and #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN240F (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.


//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN240 (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.


//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module AN241 (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;

           and #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN260F (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.


//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN310F (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN310 (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module AN311 (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;

           and #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN320F (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN320 (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module AN321 (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;

           and #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN340F (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN340 (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module AN341 (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;

           and #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN360F (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN410F (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN410 (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN420F (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN420 (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN440F (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN440 (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AN460F (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           and #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AP001 (  A );

// Verilog Port Declaration section

   input  A;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf   TI_BUF_PRIM0 ( ACC_A , A ) ;

`ifdef TI_functiononly
`else

specify


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module AP002 (  A );

// Verilog Port Declaration section

   input  A;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf   TI_BUF_PRIM0 ( ACC_A , A ) ;

`ifdef TI_functiononly
`else

specify


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF310F ( A1, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect


        and TI_AND_PRIM0  ( NODE1, B1, B2 ) ;
        nor #0 TI_NOR_PRIM0 ( Y, A1, NODE1 ) ;
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF310 ( A1, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect


        and TI_AND_PRIM0  ( NODE1, B1, B2 ) ;
        nor #0 TI_NOR_PRIM0 ( Y, A1, NODE1 ) ;
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF311F ( A1, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect

        and TI_AND_PRIM0 ( NODE1, B1, B2 ) ;
        or #0 TI_OR_PRIM0 ( Y, A1, NODE1 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF311 ( A1, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect

        and TI_AND_PRIM0 ( NODE1, B1, B2 ) ;
        or #0 TI_OR_PRIM0 ( Y, A1, NODE1 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module BF312F ( A1, B1, B2, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect

        or TI_OR_PRIM0 ( NODE1, B1, B2 ) ;
        nand #0 TI_NAND_PRIM0 ( Y, A1, NODE1 ) ;

`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module BF312 ( A1, B1, B2, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect

        or TI_OR_PRIM0 ( NODE1, B1, B2 ) ;
        nand #0 TI_NAND_PRIM0 ( Y, A1, NODE1 ) ;

`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
         
module BF313F ( A1, B1, B2, Y ) ;
     
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;

`ifdef TI_openhdl
`else
  `protect

        or TI_OR_PRIM0 ( NODE1, B1, B2 ) ;
        and #0 TI_AND_PRIM0 ( Y, A1, NODE1 ) ;

`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
         
module BF313 ( A1, B1, B2, Y ) ;
     
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;

`ifdef TI_openhdl
`else
  `protect

        or TI_OR_PRIM0 ( NODE1, B1, B2 ) ;
        and #0 TI_AND_PRIM0 ( Y, A1, NODE1 ) ;

`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF320F ( A1, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect


        and TI_AND_PRIM0  ( NODE1, B1, B2 ) ;
        nor #0 TI_NOR_PRIM0 ( Y, A1, NODE1 ) ;
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF320 ( A1, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect


        and TI_AND_PRIM0  ( NODE1, B1, B2 ) ;
        nor #0 TI_NOR_PRIM0 ( Y, A1, NODE1 ) ;
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF321F ( A1, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect

        and TI_AND_PRIM0 ( NODE1, B1, B2 ) ;
        or #0 TI_OR_PRIM0 ( Y, A1, NODE1 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF321 ( A1, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect

        and TI_AND_PRIM0 ( NODE1, B1, B2 ) ;
        or #0 TI_OR_PRIM0 ( Y, A1, NODE1 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module BF322F ( A1, B1, B2, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect

        or TI_OR_PRIM0 ( NODE1, B1, B2 ) ;
        nand #0 TI_NAND_PRIM0 ( Y, A1, NODE1 ) ;

`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module BF322 ( A1, B1, B2, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect

        or TI_OR_PRIM0 ( NODE1, B1, B2 ) ;
        nand #0 TI_NAND_PRIM0 ( Y, A1, NODE1 ) ;

`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
         
module BF323F ( A1, B1, B2, Y ) ;
     
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;

`ifdef TI_openhdl
`else
  `protect

        or TI_OR_PRIM0 ( NODE1, B1, B2 ) ;
        and #0 TI_AND_PRIM0 ( Y, A1, NODE1 ) ;

`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
         
module BF323 ( A1, B1, B2, Y ) ;
     
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;

`ifdef TI_openhdl
`else
  `protect

        or TI_OR_PRIM0 ( NODE1, B1, B2 ) ;
        and #0 TI_AND_PRIM0 ( Y, A1, NODE1 ) ;

`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF340F ( A1, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect


        and TI_AND_PRIM0  ( NODE1, B1, B2 ) ;
        nor #0 TI_NOR_PRIM0 ( Y, A1, NODE1 ) ;
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF341F ( A1, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect

        and TI_AND_PRIM0 ( NODE1, B1, B2 ) ;
        or #0 TI_OR_PRIM0 ( Y, A1, NODE1 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module BF342F ( A1, B1, B2, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect

        or TI_OR_PRIM0 ( NODE1, B1, B2 ) ;
        nand #0 TI_NAND_PRIM0 ( Y, A1, NODE1 ) ;

`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
         
module BF343F ( A1, B1, B2, Y ) ;
     
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;

`ifdef TI_openhdl
`else
  `protect

        or TI_OR_PRIM0 ( NODE1, B1, B2 ) ;
        and #0 TI_AND_PRIM0 ( Y, A1, NODE1 ) ;

`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module BF410 ( A1, A2, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


        and TI_AND_PRIM0 ( NODE1, A1, A2 ) ;
        and TI_AND_PRIM1 ( NODE2, B1, B2 ) ;
        nor #0 TI_NOR_PRIM0 ( Y, NODE1, NODE2 ) ;
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module BF411 ( A1, A2, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
        and TI_AND_PRIM0 ( NODE1, A1, A2 ) ;
        and TI_AND_PRIM1 ( NODE2, B1, B2 ) ;
        or #0 TI_OR_PRIM0 ( Y, NODE1, NODE2 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF412 ( A1, A2, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect

    // Verilog Structure section (in terms of gate prims)
        or TI_OR_PRIM0 ( NODE1, A1, A2 ) ;
        or TI_OR_PRIM1 ( NODE2, B1, B2 ) ;
        nand #0 TI_NAND_PRIM0 ( Y, NODE1, NODE2 ) ;
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF413 ( A1, A2, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        or TI_OR_PRIM0 ( NODE1, A1, A2 ) ;
        or TI_OR_PRIM1 ( NODE2, B1, B2 ) ;
        and #0 TI_AND_PRIM0 ( Y, NODE1, NODE2 ) ;
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF414 ( A1, B1, B2, B3, Y ) ;

        // Verilog Port Declaration section
       output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
        input B3 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        and TI_AND_PRIM0  ( NODE2, B1, B2, B3 ) ;
        nor #0 TI_NOR_PRIM0 ( Y, A1, NODE2 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B3 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF415 ( A1, B1, B2, B3, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
        input B3 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


        and TI_AND_PRIM0 ( NODE2, B1, B2, B3 ) ;
        or #0 TI_OR_PRIM0 ( Y, A1, NODE2 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B3 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF416 ( A1, B1, B2, B3, Y ) ;

 // Verilog Port Declaration section
       output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
        input B3 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        or  TI_OR_PRIM0 ( NODE2, B1, B2, B3 ) ;
        nand #0 TI_NAND_PRIM0 ( Y, A1, NODE2 ) ;
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B3 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF417 ( A1, B1, B2, B3, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
        input B3 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        or TI_OR_PRIM0 ( NODE2, B1, B2, B3 ) ;
        and #0 TI_AND_PRIM0 ( Y, A1, NODE2 ) ;

 `ifdef TI_functiononly
`else

       specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B3 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module BF418 ( A1, B1, C1, C2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input C1 ;
        input C2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        and TI_AND_PRIM0 ( NODE1, C1, C2 );
        or TI_OR_PRIM0 ( NODE2, B1, NODE1 ) ;
        nand #0 TI_NAND_PRIM0 ( Y, A1, NODE2 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF419 ( A1, B1, C1, C2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input C1 ;
        input C2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        and TI_AND_PRIM0 ( NODE1, C1, C2 );
        or TI_OR_PRIM0 ( NODE2, B1, NODE1 ) ;
        and #0 TI_AND_PRIM1 ( Y, A1, NODE2 ) ;
     
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF41A ( A1, B1, C1, C2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input C1 ;
        input C2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        or TI_OR_PRIM0 ( NODE1, C1, C2 );
        and TI_AND_PRIM0 ( NODE2, B1, NODE1 ) ;
        nor #0 TI_NOR_PRIM0 ( Y, A1, NODE2 ) ;
     
`ifdef TI_functiononly
`else
        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module BF41B ( A1, B1, C1, C2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input C1 ;
        input C2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


        or TI_OR_PRIM0 ( NODE1, C1, C2 );
        and TI_AND_PRIM0 ( NODE2, B1, NODE1 ) ;
        or #0 TI_OR_PRIM1 ( Y, A1, NODE2 ) ;
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module BF420 ( A1, A2, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


        and TI_AND_PRIM0 ( NODE1, A1, A2 ) ;
        and TI_AND_PRIM1 ( NODE2, B1, B2 ) ;
        nor #0 TI_NOR_PRIM0 ( Y, NODE1, NODE2 ) ;
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module BF421 ( A1, A2, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
        and TI_AND_PRIM0 ( NODE1, A1, A2 ) ;
        and TI_AND_PRIM1 ( NODE2, B1, B2 ) ;
        or #0 TI_OR_PRIM0 ( Y, NODE1, NODE2 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF422 ( A1, A2, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect

    // Verilog Structure section (in terms of gate prims)
        or TI_OR_PRIM0 ( NODE1, A1, A2 ) ;
        or TI_OR_PRIM1 ( NODE2, B1, B2 ) ;
        nand #0 TI_NAND_PRIM0 ( Y, NODE1, NODE2 ) ;
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF423 ( A1, A2, B1, B2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        or TI_OR_PRIM0 ( NODE1, A1, A2 ) ;
        or TI_OR_PRIM1 ( NODE2, B1, B2 ) ;
        and #0 TI_AND_PRIM0 ( Y, NODE1, NODE2 ) ;
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF424 ( A1, B1, B2, B3, Y ) ;

        // Verilog Port Declaration section
       output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
        input B3 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        and TI_AND_PRIM0  ( NODE2, B1, B2, B3 ) ;
        nor #0 TI_NOR_PRIM0 ( Y, A1, NODE2 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B3 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF425 ( A1, B1, B2, B3, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
        input B3 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


        and TI_AND_PRIM0 ( NODE2, B1, B2, B3 ) ;
        or #0 TI_OR_PRIM0 ( Y, A1, NODE2 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B3 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF426 ( A1, B1, B2, B3, Y ) ;

 // Verilog Port Declaration section
       output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
        input B3 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        or  TI_OR_PRIM0 ( NODE2, B1, B2, B3 ) ;
        nand #0 TI_NAND_PRIM0 ( Y, A1, NODE2 ) ;
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B3 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF427 ( A1, B1, B2, B3, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input B2 ;
        input B3 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        or TI_OR_PRIM0 ( NODE2, B1, B2, B3 ) ;
        and #0 TI_AND_PRIM0 ( Y, A1, NODE2 ) ;

 `ifdef TI_functiononly
`else

       specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B3 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module BF428 ( A1, B1, C1, C2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input C1 ;
        input C2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        and TI_AND_PRIM0 ( NODE1, C1, C2 );
        or TI_OR_PRIM0 ( NODE2, B1, NODE1 ) ;
        nand #0 TI_NAND_PRIM0 ( Y, A1, NODE2 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF429 ( A1, B1, C1, C2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input C1 ;
        input C2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        and TI_AND_PRIM0 ( NODE1, C1, C2 );
        or TI_OR_PRIM0 ( NODE2, B1, NODE1 ) ;
        and #0 TI_AND_PRIM1 ( Y, A1, NODE2 ) ;
     
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF42A ( A1, B1, C1, C2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input C1 ;
        input C2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        or TI_OR_PRIM0 ( NODE1, C1, C2 );
        and TI_AND_PRIM0 ( NODE2, B1, NODE1 ) ;
        nor #0 TI_NOR_PRIM0 ( Y, A1, NODE2 ) ;
     
`ifdef TI_functiononly
`else
        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module BF42B ( A1, B1, C1, C2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input C1 ;
        input C2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


        or TI_OR_PRIM0 ( NODE1, C1, C2 );
        and TI_AND_PRIM0 ( NODE2, B1, NODE1 ) ;
        or #0 TI_OR_PRIM1 ( Y, A1, NODE2 ) ;
`ifdef TI_functiononly
`else


        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF510 ( A1, A2, B1, B2, B3, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input B3 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


        and TI_AND_PRIM0 ( NODE1, B1, B2, B3 ) ;
        nor #0 TI_NOR_PRIM0 ( Y, NODE1, A1, A2 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B3 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF511 ( A1, A2, B1, B2, B3, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input B3 ;

    `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
     and TI_AND_PRIM0 ( NODE1, B1, B2, B3 ) ;
     or #0 TI_OR_PRIM0 ( Y, NODE1, A1, A2 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B3 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module BF512 ( A1, B1, C1, C2, C3, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input C1 ;
        input C2 ;
        input C3 ;

   `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

      or TI_OR_PRIM0 ( NODE1, C1, C2, C3 ) ;
      nand #0 TI_NAND_PRIM0 ( Y, NODE1, A1, B1 ) ;

 `ifdef TI_functiononly
`else
       specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C3 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF513 ( A1, B1, C1, C2, C3, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input C1 ;
        input C2 ;
        input C3 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


        or TI_OR_PRIM0 ( NODE1, C1, C2, C3 ) ;
        and #0 TI_AND_PRIM0 ( Y, NODE1, A1, B1 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C3 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF514 ( A1, A2, B1, B2, C1, Y ) ;

 // Verilog Port Declaration section
       output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;

  
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
      and TI_AND_PRIM0 ( NODE1, A1, A2 );
        and TI_AND_PRIM1 ( NODE2, B1, B2 );
        or TI_OR_PRIM0 ( NODE3, NODE1, NODE2 );
        nand #0 TI_NAND_PRIM0 ( Y, NODE3, C1 );
        
    `ifdef TI_functiononly
`else
    specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF515 ( A1, A2, B1, B2, C1, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        and TI_AND_PRIM0 ( NODE1, A1, A2 );
        and TI_AND_PRIM1  ( NODE2, B1, B2 );
        or TI_OR_PRIM0 ( NODE3, NODE1, NODE2 );
        and #0 TI_AND_PRIM2 ( Y, NODE3, C1 );
 `ifdef TI_functiononly
`else
       
        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module BF516 ( A1, A2, B1, B2, C1, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


        or TI_OR_PRIM0 ( NODE1, A1, A2 );
        or TI_OR_PRIM1 ( NODE2, B1, B2 );
        and  TI_AND_PRIM1 ( NODE3, NODE1, NODE2 );
        nor #0 TI_NOR_PRIM0 ( Y, NODE3, C1 );
        
 `ifdef TI_functiononly
`else
       specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF517 ( A1, A2, B1, B2, C1, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        or TI_OR_PRIM0 ( NODE1, A1, A2 );
        or TI_OR_PRIM1 ( NODE2, B1, B2 );
        and TI_AND_PRIM0 ( NODE3, NODE1, NODE2 );
        or #0 TI_OR_PRIM2 ( Y, NODE3, C1 );
        `ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF518 ( A1, A2, B1, B2, C1, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


        or TI_OR_PRIM0 ( NODE1, B1, B2 );
        and TI_AND_PRIM0 ( NODE2, NODE1, A1, A2 );
        nor #0 TI_NOR_PRIM0 ( Y, NODE2, C1 );
        
       `ifdef TI_functiononly
`else
 specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF519 ( A1, A2, B1, B2, C1, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        or TI_OR_PRIM0  ( NODE1, B1, B2 );
        and TI_AND_PRIM0 ( NODE2, NODE1, A1, A2 );
        or #0 TI_OR_PRIM1 ( Y, NODE2, C1 );
 `ifdef TI_functiononly
`else
       
        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

`endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF520 ( A1, A2, B1, B2, B3, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input B3 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


        and TI_AND_PRIM0 ( NODE1, B1, B2, B3 ) ;
        nor #0 TI_NOR_PRIM0 ( Y, NODE1, A1, A2 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B3 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF521 ( A1, A2, B1, B2, B3, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input B3 ;

    `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
     and TI_AND_PRIM0 ( NODE1, B1, B2, B3 ) ;
     or #0 TI_OR_PRIM0 ( Y, NODE1, A1, A2 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B3 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module BF522 ( A1, B1, C1, C2, C3, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input C1 ;
        input C2 ;
        input C3 ;

   `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

      or TI_OR_PRIM0 ( NODE1, C1, C2, C3 ) ;
      nand #0 TI_NAND_PRIM0 ( Y, NODE1, A1, B1 ) ;

 `ifdef TI_functiononly
`else
       specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C3 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF523 ( A1, B1, C1, C2, C3, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input B1 ;
        input C1 ;
        input C2 ;
        input C3 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


        or TI_OR_PRIM0 ( NODE1, C1, C2, C3 ) ;
        and #0 TI_AND_PRIM0 ( Y, NODE1, A1, B1 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C3 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF524 ( A1, A2, B1, B2, C1, Y ) ;

 // Verilog Port Declaration section
       output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;

  
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
      and TI_AND_PRIM0 ( NODE1, A1, A2 );
        and TI_AND_PRIM1 ( NODE2, B1, B2 );
        or TI_OR_PRIM0 ( NODE3, NODE1, NODE2 );
        nand #0 TI_NAND_PRIM0 ( Y, NODE3, C1 );
        
    `ifdef TI_functiononly
`else
    specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF525 ( A1, A2, B1, B2, C1, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        and TI_AND_PRIM0 ( NODE1, A1, A2 );
        and TI_AND_PRIM1  ( NODE2, B1, B2 );
        or TI_OR_PRIM0 ( NODE3, NODE1, NODE2 );
        and #0 TI_AND_PRIM2 ( Y, NODE3, C1 );
 `ifdef TI_functiononly
`else
       
        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module BF526 ( A1, A2, B1, B2, C1, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


        or TI_OR_PRIM0 ( NODE1, A1, A2 );
        or TI_OR_PRIM1 ( NODE2, B1, B2 );
        and  TI_AND_PRIM1 ( NODE3, NODE1, NODE2 );
        nor #0 TI_NOR_PRIM0 ( Y, NODE3, C1 );
        
 `ifdef TI_functiononly
`else
       specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF527 ( A1, A2, B1, B2, C1, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        or TI_OR_PRIM0 ( NODE1, A1, A2 );
        or TI_OR_PRIM1 ( NODE2, B1, B2 );
        and TI_AND_PRIM0 ( NODE3, NODE1, NODE2 );
        or #0 TI_OR_PRIM2 ( Y, NODE3, C1 );
        `ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF528 ( A1, A2, B1, B2, C1, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


        or TI_OR_PRIM0 ( NODE1, B1, B2 );
        and TI_AND_PRIM0 ( NODE2, NODE1, A1, A2 );
        nor #0 TI_NOR_PRIM0 ( Y, NODE2, C1 );
        
       `ifdef TI_functiononly
`else
 specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF529 ( A1, A2, B1, B2, C1, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        or TI_OR_PRIM0  ( NODE1, B1, B2 );
        and TI_AND_PRIM0 ( NODE2, NODE1, A1, A2 );
        or #0 TI_OR_PRIM1 ( Y, NODE2, C1 );
 `ifdef TI_functiononly
`else
       
        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

`endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module BF610 ( A1, A2, B1, B2, C1, C2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
        input C2 ;

 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        and TI_AND_PRIM0 ( NODE1, A1, A2 );
        and TI_AND_PRIM1 ( NODE2, B1, B2 );
        and TI_AND_PRIM2 ( NODE3, C1, C2 );
        nor #0 TI_NOR_PRIM0 ( Y, NODE1, NODE2, NODE3 ) ;

 `ifdef TI_functiononly
`else
       specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify



`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF612 ( A1, A2, B1, B2, C1, C2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
        input C2 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        or TI_OR_PRIM0 ( NODE1, A1, A2 );
        or TI_OR_PRIM1 ( NODE2, B1, B2 );
        or TI_OR_PRIM2 ( NODE3, C1, C2 );
        nand #0 TI_NAND_PRIM0 ( Y, NODE1, NODE2, NODE3 ) ;

    `ifdef TI_functiononly
`else
    specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module BF620 ( A1, A2, B1, B2, C1, C2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
        input C2 ;

 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        and TI_AND_PRIM0 ( NODE1, A1, A2 );
        and TI_AND_PRIM1 ( NODE2, B1, B2 );
        and TI_AND_PRIM2 ( NODE3, C1, C2 );
        nor #0 TI_NOR_PRIM0 ( Y, NODE1, NODE2, NODE3 ) ;

 `ifdef TI_functiononly
`else
       specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify



`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF622 ( A1, A2, B1, B2, C1, C2, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
        input C2 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        or TI_OR_PRIM0 ( NODE1, A1, A2 );
        or TI_OR_PRIM1 ( NODE2, B1, B2 );
        or TI_OR_PRIM2 ( NODE3, C1, C2 );
        nand #0 TI_NAND_PRIM0 ( Y, NODE1, NODE2, NODE3 ) ;

    `ifdef TI_functiononly
`else
    specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module BF810 ( A1, A2, B1, B2, C1, C2, D1, D2, Y ) ;

 // Verilog Port Declaration section
       output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
        input C2 ;
        input D1 ;
        input D2 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        and TI_AND_PRIM0 ( NODE1, A1, A2 );
        and TI_AND_PRIM1 ( NODE2, B1, B2 );
        and TI_AND_PRIM2 ( NODE3, C1, C2 );
        and TI_AND_PRIM3  ( NODE4, D1, D2 );
        nor #0 TI_NOR_PRIM0 ( Y, NODE1, NODE2, NODE3, NODE4 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( D1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( D2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF812 ( A1, A2, B1, B2, C1, C2, D1, D2, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
        input C2 ;
        input D1 ;
        input D2 ;

 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        or TI_OR_PRIM0 ( NODE1, A1, A2 );
        or TI_OR_PRIM1 ( NODE2, B1, B2 );
        or TI_OR_PRIM2 ( NODE3, C1, C2 );
        or TI_OR_PRIM3 ( NODE4, D1, D2 );
        nand #0 TI_NAND_PRIM0 ( Y, NODE1, NODE2, NODE3, NODE4 ) ;

   
`ifdef TI_functiononly

`else

     specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( D1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( D2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module BF820 ( A1, A2, B1, B2, C1, C2, D1, D2, Y ) ;

 // Verilog Port Declaration section
       output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
        input C2 ;
        input D1 ;
        input D2 ;
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        and TI_AND_PRIM0 ( NODE1, A1, A2 );
        and TI_AND_PRIM1 ( NODE2, B1, B2 );
        and TI_AND_PRIM2 ( NODE3, C1, C2 );
        and TI_AND_PRIM3  ( NODE4, D1, D2 );
        nor #0 TI_NOR_PRIM0 ( Y, NODE1, NODE2, NODE3, NODE4 ) ;
`ifdef TI_functiononly
`else

        specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( D1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( D2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BF822 ( A1, A2, B1, B2, C1, C2, D1, D2, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input A1 ;
        input A2 ;
        input B1 ;
        input B2 ;
        input C1 ;
        input C2 ;
        input D1 ;
        input D2 ;

 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        or TI_OR_PRIM0 ( NODE1, A1, A2 );
        or TI_OR_PRIM1 ( NODE2, B1, B2 );
        or TI_OR_PRIM2 ( NODE3, C1, C2 );
        or TI_OR_PRIM3 ( NODE4, D1, D2 );
        nand #0 TI_NAND_PRIM0 ( Y, NODE1, NODE2, NODE3, NODE4 ) ;

   
`ifdef TI_functiononly

`else

     specify
                ( A1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( A2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( B2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( C2 => Y ) = ( 0.0100, 0.0100 ) ;
                ( D1 => Y ) = ( 0.0100, 0.0100 ) ;
                ( D2 => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU110F (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU110 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU120F (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU120 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU130F (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU130 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU140F (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU140 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU150F (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU160F (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU180F (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU180 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU190F (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU190 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU1G0F (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU1G0 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU1W0 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU240 ( A, G, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A ;
        input G ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

           bufif1 #0 TI_BUFIF1_PRIM0 ( Y, A, G ) ;
`ifdef TI_functiononly
`else
       specify
                ( G => Y ) = ( 0.0100, 0.0100, 0.0100, 0.0100, 0.0100, 0.0100 ) ;
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU280 ( A, G, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A ;
        input G ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

           bufif1 #0 TI_BUFIF1_PRIM0 ( Y, A, G ) ;
`ifdef TI_functiononly
`else
       specify
                ( G => Y ) = ( 0.0100, 0.0100, 0.0100, 0.0100, 0.0100, 0.0100 ) ;
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU2G0 ( A, G, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A ;
        input G ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

           bufif1 #0 TI_BUFIF1_PRIM0 ( Y, A, G ) ;
`ifdef TI_functiononly
`else
       specify
                ( G => Y ) = ( 0.0100, 0.0100, 0.0100, 0.0100, 0.0100, 0.0100 ) ;
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module BU2P0 ( A, G, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A ;
        input G ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

           bufif1 #0 TI_BUFIF1_PRIM0 ( Y, A, G ) ;
`ifdef TI_functiononly
`else
       specify
                ( G => Y ) = ( 0.0100, 0.0100, 0.0100, 0.0100, 0.0100, 0.0100 ) ;
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2009 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

 `resetall
 `ifdef TI_verifault
      `suppress_faults
      `enable_portfaults
 `endif //TI_verifault
 
 `celldefine
 
 `ifdef TI_functiononly
     `delay_mode_distributed
     `timescale 1ps / 1ps
 `else
     `delay_mode_path
     `timescale 1ns / 1ps
 `endif //TI_functiononly
 
 // Verilog Interface section
 
 module CGN40  (CLK, EN, GCLK);
   
 // Verilog Port Declaration section
 //inputs
      input CLK ;
      input EN ;
 //outputs
      output GCLK ;
   
 `ifdef TI_verilog    
     parameter Xon = 1;
     parameter TCHKON = 1;
     wire TCHKON_NET;
     assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
 //    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
 `endif
   
 `ifdef TI_openhdl
 `else 
   `protect
      wire GVCnotifier1;
 //  Verilog Notifier declaration section
 
     reg GVCnotifier1_zd ;
 
 // Xon controlability
 
 `ifdef TI_verilog
    and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
 `endif 
 
 
       `ifdef TI_verilog
 
 // Net Declared for negative timing check
        wire  GVC_EN_EN ,  GVC_CLK_CLK  ; 
  
 
       not                 TI_INST2     (ENZ, GVC_EN_EN);
       la_nudp             TI_INST0     (ENL, ENZ, GVC_CLK_CLK, GVCnotifier1);
       or                  TI_INST3     (GCLK,ENL,GVC_CLK_CLK);
      
     `else
 
       not                 TI_INST6     (ENZ, EN);
       la_nudp             TI_INST4     (ENL, ENZ, CLK, GVCnotifier1);
       or         #0       TI_INST7     (GCLK,ENL,CLK);
   			  
      `endif//TI_verilog
   
     `ifdef TI_verilog
           cons_udp    TI_COND1  (GVC_EN_NOTEQ_ENL,ENZ , GCLK, 1'b0, 1'b1, 1'b1, 1'b1);
   
     `endif//TI_verilog
     `ifdef TI_functiononly
     
     `else
 `ifdef TI_verilog
 
     wire TCHKON_AND_GVC_EN_NOTEQ_ENL;
     and TI_AND_GVC_EN_NOTEQ_ENL (TCHKON_AND_GVC_EN_NOTEQ_ENL, GVC_EN_NOTEQ_ENL, TCHKON_NET);
 
 `endif
     
   specify    
   
     (CLK *> GCLK) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
   
         
          `ifdef TI_verilog 
          
             $setuphold(negedge CLK &&& (TCHKON_NET != 0) ,  posedge EN,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_EN_EN ); 
             $setuphold(negedge CLK &&& (TCHKON_NET != 0) ,  negedge EN,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_EN_EN ); 
             $width(posedge CLK  &&& TCHKON_AND_GVC_EN_NOTEQ_ENL != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
          
          `endif//TI_verilog
          
          
          endspecify
   
     `endif//TI_functiononly
     
     `endprotect
 `endif//TI_openhdl
 
 endmodule
 
 `endcelldefine
 
 `ifdef TI_verifault
     `nosuppress_faults
     `disable_portfaults
 `endif//TI_verifault
     
   
// Revision history:
// ----------------
//      26-Nov-2009: Mazhar, Sharavathi, Santosh. Updated #1 to #0 and updated
//                   cons_udp to have check between EN and GCLK.  Removed buf
//                   at ENL
//      27-Nov-2009: Mazhar, Sharavathi: Updated net connections so that "NOT"
//                   gate at output of latch is now placed at input of latch
//      21-Jan-2010: Mazhar. Updated to remove TI_veritime
//---------------------------------------------------------------------
// Copyright (c) 2009 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

 `resetall
 `ifdef TI_verifault
      `suppress_faults
      `enable_portfaults
 `endif //TI_verifault
 
 `celldefine
 
 `ifdef TI_functiononly
     `delay_mode_distributed
     `timescale 1ps / 1ps
 `else
     `delay_mode_path
     `timescale 1ns / 1ps
 `endif //TI_functiononly
 
 // Verilog Interface section
 
 module CGN80  (CLK, EN, GCLK);
   
 // Verilog Port Declaration section
 //inputs
      input CLK ;
      input EN ;
 //outputs
      output GCLK ;
   
 `ifdef TI_verilog    
     parameter Xon = 1;
     parameter TCHKON = 1;
     wire TCHKON_NET;
     assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
 //    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
 `endif
   
 `ifdef TI_openhdl
 `else 
   `protect
      wire GVCnotifier1;
 //  Verilog Notifier declaration section
 
     reg GVCnotifier1_zd ;
 
 // Xon controlability
 
 `ifdef TI_verilog
    and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
 `endif 
 
 
       `ifdef TI_verilog
 
 // Net Declared for negative timing check
        wire  GVC_EN_EN ,  GVC_CLK_CLK  ; 
  
 
       not                 TI_INST2     (ENZ, GVC_EN_EN);
       la_nudp             TI_INST0     (ENL, ENZ, GVC_CLK_CLK, GVCnotifier1);
       or                  TI_INST3     (GCLK,ENL,GVC_CLK_CLK);
      
     `else
 
       not                 TI_INST6     (ENZ, EN);
       la_nudp             TI_INST4     (ENL, ENZ, CLK, GVCnotifier1);
       or         #0       TI_INST7     (GCLK,ENL,CLK);
   			  
      `endif//TI_verilog
   
     `ifdef TI_verilog
           cons_udp    TI_COND1  (GVC_EN_NOTEQ_ENL,ENZ , GCLK, 1'b0, 1'b1, 1'b1, 1'b1);
   
     `endif//TI_verilog
     `ifdef TI_functiononly
     
     `else
 `ifdef TI_verilog
 
     wire TCHKON_AND_GVC_EN_NOTEQ_ENL;
     and TI_AND_GVC_EN_NOTEQ_ENL (TCHKON_AND_GVC_EN_NOTEQ_ENL, GVC_EN_NOTEQ_ENL, TCHKON_NET);
 
 `endif
     
   specify    
   
     (CLK *> GCLK) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
   
         
          `ifdef TI_verilog 
          
             $setuphold(negedge CLK &&& (TCHKON_NET != 0) ,  posedge EN,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_EN_EN ); 
             $setuphold(negedge CLK &&& (TCHKON_NET != 0) ,  negedge EN,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_EN_EN ); 
             $width(posedge CLK  &&& TCHKON_AND_GVC_EN_NOTEQ_ENL != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
          
          `endif//TI_verilog
          
          
          endspecify
   
     `endif//TI_functiononly
     
     `endprotect
 `endif//TI_openhdl
 
 endmodule
 
 `endcelldefine
 
 `ifdef TI_verifault
     `nosuppress_faults
     `disable_portfaults
 `endif//TI_verifault
     
   
// Revision history:
// ----------------
//      26-Nov-2009: Mazhar, Sharavathi, Santosh. Updated #1 to #0 and updated
//                   cons_udp to have check between EN and GCLK.  Removed buf
//                   at ENL
//      27-Nov-2009: Mazhar, Sharavathi: Updated net connections so that "NOT"
//                   gate at output of latch is now placed at input of latch
//      21-Jan-2010: Mazhar. Updated to remove TI_veritime
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

 `resetall
 `ifdef TI_verifault
      `suppress_faults
      `enable_portfaults
 `endif //TI_verifault
 
 `celldefine
 
 `ifdef TI_functiononly
     `delay_mode_distributed
     `timescale 1ps/1ps
 `else
     `delay_mode_path
     `timescale 1ns / 1ps
 `endif //TI_functiononly
 
 // Verilog Interface section
 
 module CGNT40 (CLK, EN, TE, GCLK);
  
 // Verilog Port Declaration section
 //inputs
      input CLK ;
      input EN ;
      input TE ;
 //outputs
      output GCLK ;
   
   
 `ifdef TI_verilog    
     parameter Xon = 1;
     parameter TCHKON = 1;
     wire TCHKON_NET;
     assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
 //    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
 `endif
   
 `ifdef TI_openhdl
 `else 
   `protect
      wire GVCnotifier1;
 //  Verilog Notifier declaration section
 
     reg GVCnotifier1_zd ;
 
 // Xon controlability
 
 `ifdef TI_verilog
    and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
 `endif 
 
 
       `ifdef TI_verilog
 
 // Net Declared for negative timing check
      wire GVC_EN_EN , GVC_CLK_CLK , GVC_TE_TE ;
   
       nor                 TI_INST4     (D_INT_inv, GVC_EN_EN, GVC_TE_TE); 
       la_nudp             TI_INST0     (ENL, D_INT_inv, GVC_CLK_CLK, GVCnotifier1);
       or                  TI_INST3     (GCLK,ENL,GVC_CLK_CLK);
      
     `else
       nor                 TI_INST4     (D_INT_inv, EN, TE); 
       la_nudp             TI_INST0     (ENL, D_INT_inv, CLK, GVCnotifier1);
       or        #0        TI_INST3     (GCLK,ENL,CLK);
   
   
      `endif//TI_verilog
   
     `ifdef TI_verilog
       cons_udp            TI_COND0     (GVC_EN_NOTEQ_ENL, D_INT_inv, GCLK, 1'b0, 1'b1, 1'b1, 1'b1);
   
     `endif//TI_verilog
 
     `ifdef TI_functiononly
     
     `else
 `ifdef TI_verilog
     wire TCHKON_AND_GVC_EN_NOTEQ_ENL;
 
     not TI_COND2 (EN_inv, GVC_EN_EN);
     not TI_COND3 (TE_inv, GVC_TE_TE);
 
     and TI_COND4 (TCHKON_AND_EN_inv, EN_inv, TCHKON_NET);
     and TI_COND5 (TCHKON_AND_TE_inv, TE_inv, TCHKON_NET);
 
     and TI_AND_GVC_EN_NOTEQ_ENL (TCHKON_AND_GVC_EN_NOTEQ_ENL, GVC_EN_NOTEQ_ENL, TCHKON_NET);
 
 `endif
     
   specify    
   
     (CLK *> GCLK) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
   
          
          `ifdef TI_verilog 
          
             $setuphold(negedge CLK ,  posedge EN,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_TE_inv != 0, GVC_CLK_CLK, GVC_EN_EN ); 
             $setuphold(negedge CLK ,  negedge EN,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_TE_inv != 0, GVC_CLK_CLK, GVC_EN_EN ); 
             $setuphold(negedge CLK ,  posedge TE,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_EN_inv != 0, GVC_CLK_CLK, GVC_TE_TE ); 
             $setuphold(negedge CLK ,  negedge TE,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_EN_inv != 0, GVC_CLK_CLK, GVC_TE_TE ); 
             $width(posedge CLK  &&& TCHKON_AND_GVC_EN_NOTEQ_ENL != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
          
          `endif//TI_verilog
          
          
          endspecify
   
     `endif//TI_functiononly
     
     `endprotect
 `endif//TI_openhdl
 
 endmodule
 
 `endcelldefine
 
 `ifdef TI_verifault
     `nosuppress_faults
     `disable_portfaults
 `endif//TI_verifault


// Revision history:
// ----------------
//      26-Nov-2009: Mazhar, Sharavathi, Santosh. Updated #1 to #0 and updated
//                   cons_udp to have check between EN and GCLK.  Removed buf
//                   at ENL
//      27-Nov-2009: Mazhar, Sharavathi: Updated net connections to be similar
//                   to that in asic models (i.e., "NOT" gate at output of 
//                   latch is now placed at input of latch
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

 `resetall
 `ifdef TI_verifault
      `suppress_faults
      `enable_portfaults
 `endif //TI_verifault
 
 `celldefine
 
 `ifdef TI_functiononly
     `delay_mode_distributed
     `timescale 1ps/1ps
 `else
     `delay_mode_path
     `timescale 1ns / 1ps
 `endif //TI_functiononly
 
 // Verilog Interface section
 
 module CGNT80 (CLK, EN, TE, GCLK);
  
 // Verilog Port Declaration section
 //inputs
      input CLK ;
      input EN ;
      input TE ;
 //outputs
      output GCLK ;
   
   
 `ifdef TI_verilog    
     parameter Xon = 1;
     parameter TCHKON = 1;
     wire TCHKON_NET;
     assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
 //    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
 `endif
   
 `ifdef TI_openhdl
 `else 
   `protect
      wire GVCnotifier1;
 //  Verilog Notifier declaration section
 
     reg GVCnotifier1_zd ;
 
 // Xon controlability
 
 `ifdef TI_verilog
    and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
 `endif 
 
 
       `ifdef TI_verilog
 
 // Net Declared for negative timing check
      wire GVC_EN_EN , GVC_CLK_CLK , GVC_TE_TE ;
   
       nor                 TI_INST4     (D_INT_inv, GVC_EN_EN, GVC_TE_TE); 
       la_nudp             TI_INST0     (ENL, D_INT_inv, GVC_CLK_CLK, GVCnotifier1);
       or                  TI_INST3     (GCLK,ENL,GVC_CLK_CLK);
      
     `else
       nor                 TI_INST4     (D_INT_inv, EN, TE); 
       la_nudp             TI_INST0     (ENL, D_INT_inv, CLK, GVCnotifier1);
       or        #0        TI_INST3     (GCLK,ENL,CLK);
   
   
      `endif//TI_verilog
   
     `ifdef TI_verilog
       cons_udp            TI_COND0     (GVC_EN_NOTEQ_ENL, D_INT_inv, GCLK, 1'b0, 1'b1, 1'b1, 1'b1);
   
     `endif//TI_verilog
 
     `ifdef TI_functiononly
     
     `else
 `ifdef TI_verilog
     wire TCHKON_AND_GVC_EN_NOTEQ_ENL;
 
     not TI_COND2 (EN_inv, GVC_EN_EN);
     not TI_COND3 (TE_inv, GVC_TE_TE);
 
     and TI_COND4 (TCHKON_AND_EN_inv, EN_inv, TCHKON_NET);
     and TI_COND5 (TCHKON_AND_TE_inv, TE_inv, TCHKON_NET);
 
     and TI_AND_GVC_EN_NOTEQ_ENL (TCHKON_AND_GVC_EN_NOTEQ_ENL, GVC_EN_NOTEQ_ENL, TCHKON_NET);
 
 `endif
     
   specify    
   
     (CLK *> GCLK) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
   
          
          `ifdef TI_verilog 
          
             $setuphold(negedge CLK ,  posedge EN,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_TE_inv != 0, GVC_CLK_CLK, GVC_EN_EN ); 
             $setuphold(negedge CLK ,  negedge EN,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_TE_inv != 0, GVC_CLK_CLK, GVC_EN_EN ); 
             $setuphold(negedge CLK ,  posedge TE,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_EN_inv != 0, GVC_CLK_CLK, GVC_TE_TE ); 
             $setuphold(negedge CLK ,  negedge TE,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_EN_inv != 0, GVC_CLK_CLK, GVC_TE_TE ); 
             $width(posedge CLK  &&& TCHKON_AND_GVC_EN_NOTEQ_ENL != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
          
          `endif//TI_verilog
          
          
          endspecify
   
     `endif//TI_functiononly
     
     `endprotect
 `endif//TI_openhdl
 
 endmodule
 
 `endcelldefine
 
 `ifdef TI_verifault
     `nosuppress_faults
     `disable_portfaults
 `endif//TI_verifault


// Revision history:
// ----------------
//      26-Nov-2009: Mazhar, Sharavathi, Santosh. Updated #1 to #0 and updated
//                   cons_udp to have check between EN and GCLK.  Removed buf
//                   at ENL
//      27-Nov-2009: Mazhar, Sharavathi: Updated net connections to be similar
//                   to that in asic models (i.e., "NOT" gate at output of 
//                   latch is now placed at input of latch
//---------------------------------------------------------------------
// Copyright (c) 2009 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

 `resetall
 `ifdef TI_verifault
      `suppress_faults
      `enable_portfaults
 `endif //TI_verifault
 
 `celldefine
 
 `ifdef TI_functiononly
     `delay_mode_distributed
     `timescale 1ps / 1ps
 `else
     `delay_mode_path
     `timescale 1ns / 1ps
 `endif //TI_functiononly
 
 // Verilog Interface section
 
 module CGP40 (CLK, EN, GCLK);
   
 // Verilog Port Declaration section
 //inputs
      input CLK ;
      input EN ;
 //outputs
      output GCLK ;
   
 `ifdef TI_verilog    
     parameter Xon = 1;
     parameter TCHKON = 1;
     wire TCHKON_NET;
     assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
 //    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
 `endif
   
 `ifdef TI_openhdl
 `else 
   `protect
      wire GVCnotifier1;
 //  Verilog Notifier declaration section
 
     reg GVCnotifier1_zd ;
 
 // Xon controlability
 
 `ifdef TI_verilog
    and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
 `endif 
 
 
       `ifdef TI_verilog
 
 // Net Declared for negative timing check
 
          wire GVC_CLK_CLK , GVC_EN_EN ;
   
   
         not                 TI_INST0     (IINVnet1, GVC_CLK_CLK);
         la_nudp             TI_INST1     (ENL, GVC_EN_EN, IINVnet1, GVCnotifier1);
         and                 TI_INST4     (GCLK,ENL,GVC_CLK_CLK);
    
     `else
           
          not                 TI_INST7     (IINVnet1, CLK);
          la_nudp             TI_INST8     (ENL, EN, IINVnet1, GVCnotifier1);
          and     #0          TI_INST10     (GCLK,ENL,CLK);
 
      `endif//TI_verilog
   
     `ifdef TI_verilog
     
        //  Logic enabling constraint check statements for verilog/verifault
         cons_udp            TI_COND1     (GVC_EN_NOTEQ_ENL, GVC_EN_EN, GCLK, 1'b0, 1'b1, 1'b1, 1'b1);
               
     `endif//TI_verilog
     `ifdef TI_functiononly
     
     `else
 `ifdef TI_verilog
 
     wire TCHKON_AND_GVC_EN_NOTEQ_ENL;
     and TI_AND_GVC_EN_NOTEQ_ENL (TCHKON_AND_GVC_EN_NOTEQ_ENL, GVC_EN_NOTEQ_ENL, TCHKON_NET);
 
 `endif
     
   
   specify    
   
     (CLK *> GCLK) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);  
   
          
          `ifdef TI_verilog 
          
             $setuphold(posedge CLK &&& (TCHKON_NET != 0) ,  posedge EN,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_EN_EN ); 
             $setuphold(posedge CLK &&& (TCHKON_NET != 0) ,  negedge EN,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_EN_EN ); 
             $width(negedge CLK  &&& TCHKON_AND_GVC_EN_NOTEQ_ENL != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
          
          `endif//TI_verilog
          
          
          endspecify
     `endif//TI_functiononly
     
     `endprotect
 `endif//TI_openhdl
 
 endmodule
 
 `endcelldefine
 
 `ifdef TI_verifault
     `nosuppress_faults
     `disable_portfaults
 `endif//TI_verifault
     
  
// Revision history:
// ----------------
//      26-Nov-2009: Mazhar, Sharavathi, Santosh. Updated #1 to #0 and updated
//                   cons_udp to have check between EN and GCLK.  Removed buf
//                   at ENL
//      21-Jan-2010: Mazhar. Updated to remove TI_veritime
//---------------------------------------------------------------------
// Copyright (c) 2009 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

 `resetall
 `ifdef TI_verifault
      `suppress_faults
      `enable_portfaults
 `endif //TI_verifault
 
 `celldefine
 
 `ifdef TI_functiononly
     `delay_mode_distributed
     `timescale 1ps / 1ps
 `else
     `delay_mode_path
     `timescale 1ns / 1ps
 `endif //TI_functiononly
 
 // Verilog Interface section
 
 module CGP80 (CLK, EN, GCLK);
   
 // Verilog Port Declaration section
 //inputs
      input CLK ;
      input EN ;
 //outputs
      output GCLK ;
   
 `ifdef TI_verilog    
     parameter Xon = 1;
     parameter TCHKON = 1;
     wire TCHKON_NET;
     assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
 //    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
 `endif
   
 `ifdef TI_openhdl
 `else 
   `protect
      wire GVCnotifier1;
 //  Verilog Notifier declaration section
 
     reg GVCnotifier1_zd ;
 
 // Xon controlability
 
 `ifdef TI_verilog
    and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
 `endif 
 
 
       `ifdef TI_verilog
 
 // Net Declared for negative timing check
 
          wire GVC_CLK_CLK , GVC_EN_EN ;
   
   
         not                 TI_INST0     (IINVnet1, GVC_CLK_CLK);
         la_nudp             TI_INST1     (ENL, GVC_EN_EN, IINVnet1, GVCnotifier1);
         and                 TI_INST4     (GCLK,ENL,GVC_CLK_CLK);
    
     `else
           
          not                 TI_INST7     (IINVnet1, CLK);
          la_nudp             TI_INST8     (ENL, EN, IINVnet1, GVCnotifier1);
          and     #0          TI_INST10     (GCLK,ENL,CLK);
 
      `endif//TI_verilog
   
     `ifdef TI_verilog
     
        //  Logic enabling constraint check statements for verilog/verifault
         cons_udp            TI_COND1     (GVC_EN_NOTEQ_ENL, GVC_EN_EN, GCLK, 1'b0, 1'b1, 1'b1, 1'b1);
               
     `endif//TI_verilog
     `ifdef TI_functiononly
     
     `else
 `ifdef TI_verilog
 
     wire TCHKON_AND_GVC_EN_NOTEQ_ENL;
     and TI_AND_GVC_EN_NOTEQ_ENL (TCHKON_AND_GVC_EN_NOTEQ_ENL, GVC_EN_NOTEQ_ENL, TCHKON_NET);
 
 `endif
     
   
   specify    
   
     (CLK *> GCLK) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);  
   
          
          `ifdef TI_verilog 
          
             $setuphold(posedge CLK &&& (TCHKON_NET != 0) ,  posedge EN,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_EN_EN ); 
             $setuphold(posedge CLK &&& (TCHKON_NET != 0) ,  negedge EN,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_EN_EN ); 
             $width(negedge CLK  &&& TCHKON_AND_GVC_EN_NOTEQ_ENL != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
          
          `endif//TI_verilog
          
          
          endspecify
     `endif//TI_functiononly
     
     `endprotect
 `endif//TI_openhdl
 
 endmodule
 
 `endcelldefine
 
 `ifdef TI_verifault
     `nosuppress_faults
     `disable_portfaults
 `endif//TI_verifault
     
  
// Revision history:
// ----------------
//      26-Nov-2009: Mazhar, Sharavathi, Santosh. Updated #1 to #0 and updated
//                   cons_udp to have check between EN and GCLK.  Removed buf
//                   at ENL
//      21-Jan-2010: Mazhar. Updated to remove TI_veritime
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
     `suppress_faults
     `enable_portfaults
`endif //TI_verifault

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
     `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif //TI_functiononly

// Verilog Interface section

module CGPT40 (CLK, EN, TE, GCLK);
 
// Verilog Port Declaration section
//inputs
     input CLK ;
     input EN ;
     input TE ;
//outputs
     output GCLK ;
  
`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif
  
`ifdef TI_openhdl
`else 
  `protect
     wire GVCnotifier1;
//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
`endif 


      `ifdef TI_verilog

// Net Declared for negative timing check

         wire GVC_CLK_CLK , GVC_EN_EN , GVC_TE_TE;
  
         or                  TI_INST5     (D_INT, GVC_EN_EN, GVC_TE_TE); 
         not                 TI_INST0     (IINVnet1, GVC_CLK_CLK);
         la_nudp             TI_INST1     (ENL, D_INT, IINVnet1, GVCnotifier1);
         and                 TI_INST4     (GCLK,ENL,GVC_CLK_CLK);

      `else
          
         or                  TI_INST6     (D_INT, EN, TE); 
         not                 TI_INST7     (IINVnet1, CLK);
         la_nudp             TI_INST8     (ENL, D_INT, IINVnet1, GVCnotifier1);
         and        #0       TI_INST10     (GCLK,ENL,CLK);


     `endif//TI_verilog
  
    `ifdef TI_verilog
    
       //  Logic enabling constraint check statements for verilog/verifault
         cons_udp            TI_COND0     (GVC_EN_NOTEQ_ENL, D_INT, GCLK, 1'b0, 1'b1, 1'b1, 1'b1);
              
    `endif//TI_verilog

    `ifdef TI_functiononly
    
     `else
`ifdef TI_verilog

 wire TCHKON_AND_GVC_EN_NOTEQ_ENL;

    not TI_COND2 (EN_inv, GVC_EN_EN);
    not TI_COND3 (TE_inv, GVC_TE_TE);

    and TI_COND4 (TCHKON_AND_EN_inv, EN_inv, TCHKON_NET);
    and TI_COND5 (TCHKON_AND_TE_inv, TE_inv, TCHKON_NET);

 and TI_AND_GVC_EN_NOTEQ_ENL (TCHKON_AND_GVC_EN_NOTEQ_ENL, GVC_EN_NOTEQ_ENL, TCHKON_NET);

`endif
    
         specify
           
             ( CLK *> GCLK) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
         
         
         `ifdef TI_verilog 
         
            $setuphold(posedge CLK ,  posedge EN,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_TE_inv != 0, GVC_CLK_CLK, GVC_EN_EN ); 
            $setuphold(posedge CLK ,  negedge EN,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_TE_inv != 0, GVC_CLK_CLK, GVC_EN_EN ); 
            $setuphold(posedge CLK ,  posedge TE,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_EN_inv != 0, GVC_CLK_CLK, GVC_TE_TE ); 
            $setuphold(posedge CLK ,  negedge TE,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_EN_inv != 0, GVC_CLK_CLK, GVC_TE_TE ); 
            $width(negedge CLK  &&& TCHKON_AND_GVC_EN_NOTEQ_ENL != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
         
         `endif//TI_verilog
         
         
         endspecify
    `endif//TI_functiononly
    
    `endprotect
`endif//TI_openhdl

endmodule

`endcelldefine

`ifdef TI_verifault
    `nosuppress_faults
    `disable_portfaults
`endif//TI_verifault
    
// Revision history:
// ----------------
//      26-Nov-2009: Mazhar, Sharavathi, Santosh. Updated #1 to #0 and updated
//                   cons_udp to have check between EN and GCLK.  Removed buf
//                   at ENL
// v1.2 12-Sep-2007 :Dundappa.
//                   Added the default delay of 1 for the output pins.
// v1.1	 11-Jan-2006 removed "TI_veritime" defination from models
// v1.0  10-Jan-2006 Currently the model is flagging setup/hold violation between CLK and TE pins
//                   and setup/hold vilation between CLK  and EN pins irrespective of the
//                   EN or TE pins respectively.
//                   This is not correct as EN is ORed with TE So if any one signal is high
//                   The other pin should not be checked for setup/hold timings against CLK pin
//                   TCHKON_AND_TE_inv != 0 and TCHKON_AND_EN_inv != 0"  is used
//                   to check the status of other pin before checking the setup/hold violations.
//                   Updated for "TCHKON_AND_TE_inv != 0" and 
//		     removed "TI_veritime" from models
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
     `suppress_faults
     `enable_portfaults
`endif //TI_verifault

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
     `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif //TI_functiononly

// Verilog Interface section

module CGPT80 (CLK, EN, TE, GCLK);
 
// Verilog Port Declaration section
//inputs
     input CLK ;
     input EN ;
     input TE ;
//outputs
     output GCLK ;
  
`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif
  
`ifdef TI_openhdl
`else 
  `protect
     wire GVCnotifier1;
//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
`endif 


      `ifdef TI_verilog

// Net Declared for negative timing check

         wire GVC_CLK_CLK , GVC_EN_EN , GVC_TE_TE;
  
         or                  TI_INST5     (D_INT, GVC_EN_EN, GVC_TE_TE); 
         not                 TI_INST0     (IINVnet1, GVC_CLK_CLK);
         la_nudp             TI_INST1     (ENL, D_INT, IINVnet1, GVCnotifier1);
         and                 TI_INST4     (GCLK,ENL,GVC_CLK_CLK);

      `else
          
         or                  TI_INST6     (D_INT, EN, TE); 
         not                 TI_INST7     (IINVnet1, CLK);
         la_nudp             TI_INST8     (ENL, D_INT, IINVnet1, GVCnotifier1);
         and        #0       TI_INST10     (GCLK,ENL,CLK);


     `endif//TI_verilog
  
    `ifdef TI_verilog
    
       //  Logic enabling constraint check statements for verilog/verifault
         cons_udp            TI_COND0     (GVC_EN_NOTEQ_ENL, D_INT, GCLK, 1'b0, 1'b1, 1'b1, 1'b1);
              
    `endif//TI_verilog

    `ifdef TI_functiononly
    
     `else
`ifdef TI_verilog

 wire TCHKON_AND_GVC_EN_NOTEQ_ENL;

    not TI_COND2 (EN_inv, GVC_EN_EN);
    not TI_COND3 (TE_inv, GVC_TE_TE);

    and TI_COND4 (TCHKON_AND_EN_inv, EN_inv, TCHKON_NET);
    and TI_COND5 (TCHKON_AND_TE_inv, TE_inv, TCHKON_NET);

 and TI_AND_GVC_EN_NOTEQ_ENL (TCHKON_AND_GVC_EN_NOTEQ_ENL, GVC_EN_NOTEQ_ENL, TCHKON_NET);

`endif
    
         specify
           
             ( CLK *> GCLK) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
         
         
         `ifdef TI_verilog 
         
            $setuphold(posedge CLK ,  posedge EN,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_TE_inv != 0, GVC_CLK_CLK, GVC_EN_EN ); 
            $setuphold(posedge CLK ,  negedge EN,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_TE_inv != 0, GVC_CLK_CLK, GVC_EN_EN ); 
            $setuphold(posedge CLK ,  posedge TE,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_EN_inv != 0, GVC_CLK_CLK, GVC_TE_TE ); 
            $setuphold(posedge CLK ,  negedge TE,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_EN_inv != 0, GVC_CLK_CLK, GVC_TE_TE ); 
            $width(negedge CLK  &&& TCHKON_AND_GVC_EN_NOTEQ_ENL != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
         
         `endif//TI_verilog
         
         
         endspecify
    `endif//TI_functiononly
    
    `endprotect
`endif//TI_openhdl

endmodule

`endcelldefine

`ifdef TI_verifault
    `nosuppress_faults
    `disable_portfaults
`endif//TI_verifault
    
// Revision history:
// ----------------
//      26-Nov-2009: Mazhar, Sharavathi, Santosh. Updated #1 to #0 and updated
//                   cons_udp to have check between EN and GCLK.  Removed buf
//                   at ENL
// v1.2 12-Sep-2007 :Dundappa.
//                   Added the default delay of 1 for the output pins.
// v1.1	 11-Jan-2006 removed "TI_veritime" defination from models
// v1.0  10-Jan-2006 Currently the model is flagging setup/hold violation between CLK and TE pins
//                   and setup/hold vilation between CLK  and EN pins irrespective of the
//                   EN or TE pins respectively.
//                   This is not correct as EN is ORed with TE So if any one signal is high
//                   The other pin should not be checked for setup/hold timings against CLK pin
//                   TCHKON_AND_TE_inv != 0 and TCHKON_AND_EN_inv != 0"  is used
//                   to check the status of other pin before checking the setup/hold violations.
//                   Updated for "TCHKON_AND_TE_inv != 0" and 
//		     removed "TI_veritime" from models
//---------------------------------------------------------------------
// Copyright (c) 2002 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

`resetall

`ifdef TI_functiononly
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

primitive cons_udp
`protect
(out, in1, in2, in3, clk, clrz, prez);
   input  in1, in2, in3, clk, clrz, prez;
   output out; 
   table   
// in1   in2   in3   clk   clrz prez : out
   ?     ?     ?     ?     0    ?    : 0 ; // active clrz
   ?     ?     ?     ?     ?    0    : 0 ; // active prez

   0     ?     0     0     1    1    : 0 ; // in1 == in3 ; clk == 0
   1     ?     1     0     1    1    : 0 ; //    "
   x     ?     x     0     1    1    : 0 ; //    "

   0     ?     0     0     x    1    : 0 ; // in1 == in3 ; clk == 0
   1     ?     1     0     1    x    : 0 ; //    "

   0     0     ?     1     1    1    : 0 ; // in1 == in2 ; clk == 1
   1     1     ?     1     1    1    : 0 ; //    "
   x     x     ?     1     1    1    : 0 ; //    "

   0     0     ?     1     x    1    : 0 ; // in1 == in2 ; clk == 1 ; clrz = x;
   1     1     ?     1     x    1    : 0 ; //    "
   x     x     ?     1     x    1    : 0 ; //    "

   0     0     ?     1     1    x    : 0 ; // in1 == in2 ; clk == 1 ; prez = x;
   1     1     ?     1     1    x    : 0 ; //    "
   x     x     ?     1     1    x    : 0 ; //    "

   0     0     0     x     1    1    : 0 ; // in1 == in2 == in3 ; clk = x
   1     1     1     x     1    1    : 0 ; //    "
   x     x     x     x     1    1    : 0 ; //    "

   0     0     0     x     x    1    : 0 ; //    "     ; clk == x
   1     1     1     x     1    x    : 0 ; //    "     ; clk == x

   1     1     1     x     x    1    : 0 ; // clrz = x ; clk == x
   1     1     1     x     x    x    : 0 ; // clrz=x,prez=x ; clk == x
   endtable
`endprotect
endprimitive 

// Revision history:
// ----------------
// v1.2  08-Jun-1999  Changing 10ps to 1ps
// v1.1  17-Mar-1999 24 date and time created 99/03/17 17
// 19 Dec 2006 : Sharavathi : changed the timescale for functiononly option to 
//                            1ns/1ps
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module CTB15 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module CTB20 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module CTB25 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module CTB30 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module CTB35 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module CTB40 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module CTB45 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module CTB50 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module CTB55 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module CTB60 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module CTB65 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module CTB70 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module CTI15 ( A, Y ) ;
// Verilog Port Declaration section

        input A ;
        output Y ;
	
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not #0 TI_NOT_PRIM0( Y, A ) ;
	
`ifdef TI_functiononly
`else

        specify
                ( A -=> Y ) =  0.01 ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 11-Sep-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.
//v1.0 19 Apr 2006 : Shara : modified the timing path to have
//                       -=> instead of "*>" 

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module CTI20 ( A, Y ) ;
// Verilog Port Declaration section

        input A ;
        output Y ;
	
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not #0 TI_NOT_PRIM0( Y, A ) ;
	
`ifdef TI_functiononly
`else

        specify
                ( A -=> Y ) =  0.01 ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 11-Sep-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.
//v1.0 19 Apr 2006 : Shara : modified the timing path to have
//                       -=> instead of "*>" 

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module CTI25 ( A, Y ) ;
// Verilog Port Declaration section

        input A ;
        output Y ;
	
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not #0 TI_NOT_PRIM0( Y, A ) ;
	
`ifdef TI_functiononly
`else

        specify
                ( A -=> Y ) =  0.01 ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 11-Sep-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.
//v1.0 19 Apr 2006 : Shara : modified the timing path to have
//                       -=> instead of "*>" 

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module CTI30 ( A, Y ) ;
// Verilog Port Declaration section

        input A ;
        output Y ;
	
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not #0 TI_NOT_PRIM0( Y, A ) ;
	
`ifdef TI_functiononly
`else

        specify
                ( A -=> Y ) =  0.01 ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 11-Sep-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.
//v1.0 19 Apr 2006 : Shara : modified the timing path to have
//                       -=> instead of "*>" 

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module CTI35 ( A, Y ) ;
// Verilog Port Declaration section

        input A ;
        output Y ;
	
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not #0 TI_NOT_PRIM0( Y, A ) ;
	
`ifdef TI_functiononly
`else

        specify
                ( A -=> Y ) =  0.01 ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 11-Sep-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.
//v1.0 19 Apr 2006 : Shara : modified the timing path to have
//                       -=> instead of "*>" 

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module CTI40 ( A, Y ) ;
// Verilog Port Declaration section

        input A ;
        output Y ;
	
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not #0 TI_NOT_PRIM0( Y, A ) ;
	
`ifdef TI_functiononly
`else

        specify
                ( A -=> Y ) =  0.01 ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 11-Sep-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.
//v1.0 19 Apr 2006 : Shara : modified the timing path to have
//                       -=> instead of "*>" 

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module CTI45 ( A, Y ) ;
// Verilog Port Declaration section

        input A ;
        output Y ;
	
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not #0 TI_NOT_PRIM0( Y, A ) ;
	
`ifdef TI_functiononly
`else

        specify
                ( A -=> Y ) =  0.01 ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 11-Sep-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.
//v1.0 19 Apr 2006 : Shara : modified the timing path to have
//                       -=> instead of "*>" 

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module CTI50 ( A, Y ) ;
// Verilog Port Declaration section

        input A ;
        output Y ;
	
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not #0 TI_NOT_PRIM0( Y, A ) ;
	
`ifdef TI_functiononly
`else

        specify
                ( A -=> Y ) =  0.01 ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 11-Sep-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.
//v1.0 19 Apr 2006 : Shara : modified the timing path to have
//                       -=> instead of "*>" 

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module CTI55 ( A, Y ) ;
// Verilog Port Declaration section

        input A ;
        output Y ;
	
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not #0 TI_NOT_PRIM0( Y, A ) ;
	
`ifdef TI_functiononly
`else

        specify
                ( A -=> Y ) =  0.01 ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 11-Sep-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.
//v1.0 19 Apr 2006 : Shara : modified the timing path to have
//                       -=> instead of "*>" 

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module CTI60 ( A, Y ) ;
// Verilog Port Declaration section

        input A ;
        output Y ;
	
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not #0 TI_NOT_PRIM0( Y, A ) ;
	
`ifdef TI_functiononly
`else

        specify
                ( A -=> Y ) =  0.01 ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 11-Sep-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.
//v1.0 19 Apr 2006 : Shara : modified the timing path to have
//                       -=> instead of "*>" 

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module CTI65 ( A, Y ) ;
// Verilog Port Declaration section

        input A ;
        output Y ;
	
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not #0 TI_NOT_PRIM0( Y, A ) ;
	
`ifdef TI_functiononly
`else

        specify
                ( A -=> Y ) =  0.01 ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 11-Sep-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.
//v1.0 19 Apr 2006 : Shara : modified the timing path to have
//                       -=> instead of "*>" 

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section
module CTI70 ( A, Y ) ;
// Verilog Port Declaration section

        input A ;
        output Y ;
	
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not #0 TI_NOT_PRIM0( Y, A ) ;
	
`ifdef TI_functiononly
`else

        specify
                ( A -=> Y ) =  0.01 ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 11-Sep-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.
//v1.0 19 Apr 2006 : Shara : modified the timing path to have
//                       -=> instead of "*>" 

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2002 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

`resetall
`ifdef TI_functiononly
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif
primitive dffqzudp
`protect
(qz, clrz, prez, q);
input clrz, prez, q;
output qz;
   table
//    clrz prez  q  :  qz
       ?    0    ?  :  0;
       0    1    ?  :  1;
       ?    1    0  :  1;
       1    ?    1  :  0;
   endtable
`endprotect
endprimitive 


// Revision history:
// ----------------
// v1.2  08-Jun-1999  Changing 10ps to 1ps
// v1.1  17-Mar-1999 24 date and time created 99/03/17 17
// v1.2  08-Jun-1999  Changing 10ps to 1ps
// v1.1  17-Mar-1999 24 date and time created 99/03/17 17
// v1.2  08-Jun-1999  Changing 10ps to 1ps
// v1.1  17-Mar-1999 24 date and time created 99/03/17 17
// 19 Dec 2006 : Sharavathi : changed the timescale for functiononly option to 
//                            1ns/1ps
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2002 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

`resetall
`ifdef TI_functiononly
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif
primitive dlaudp(q, d, c, clr, pre, nt);

input d, c, clr, pre, nt;
output q;
reg q;

table
//  d   c   clr   pre   nt  : q :  q;
    *   ?    1     0    ?   : ? :  1;
    ?   *    1     0    ?   : ? :  1;
    ?   ?   (?1)   0    ?   : ? :  1;
    ?   ?    1    (?0)  ?   : ? :  1;

    *   ?    0     0    ?   : ? :  0;
    ?   *    0     0    ?   : ? :  0;
    ?   ?   (?0)   0    ?   : ? :  0;
    ?   ?    0    (?0)  ?   : ? :  0;

    ?   ?   (?0)   1    ?   : ? :  0;
    *   ?    0     1    ?   : ? :  0;
    ?   *    0     1    ?   : ? :  0;
    ?   ?    0    (?1)  ?   : ? :  0;
 
   (?1) ?    1     ?    ?   : 1 :  1;
    1   ?   (?1)   ?    ?   : 1 :  1;
    1   ?    1     *    ?   : 1 :  1;
    1   *    1     ?    ?   : 1 :  1;

   (?0) ?    ?     1    ?   : 0 :  0;
    0   ?    ?    (?1)  ?   : 0 :  0;
    0   *    ?     1    ?   : 0 :  0;
    0   ?    *     1    ?   : 0 :  0;

    ?  (?0)  1     1    ?   : ? :  -;
    ?   0   (?1)   1    ?   : ? :  -;
    ?   0    1    (?1)  ?   : ? :  -;
    *   0    1     1    ?   : ? :  -;

//reduction of pessimism

   (?0) 1    ?     1    ?   : ? :  0;
    0  (?1)  ?     1    ?   : ? :  0;
    0   1    ?    (?1)  ?   : ? :  0;
    0   1    *     1    ?   : ? :  0;

   (?1) 1    1     ?    ?   : ? :  1;
    1  (?1)  1     ?    ?   : ? :  1;
    1   1   (?1)   ?    ?   : ? :  1;
    1   1    1     *    ?   : ? :  1;

    ?  (?0)  x     1    ?   : 0 :  0;
    ?   0   (?x)   1    ?   : 0 :  0;
    ?   0    x    (?1)  ?   : 0 :  0;
    *   0    x     1    ?   : 0 :  0;

    ?  (?0)  1     x    ?   : 1 :  1;
    ?   0   (?1)   x    ?   : 1 :  1;
    ?   0    1    (?x)  ?   : 1 :  1;
    *   0    1     x    ?   : 1 :  1; 

    *   ?    0     x    ?   : ? :  0; 
    ?   *    0     x    ?   : ? :  0; 
    ?   ?   (?0)   x    ?   : ? :  0; 
    ?   ?    0    (?x)  ?   : ? :  0; 

    ?   ?    ?     ?    *   : ? :  x;

endtable
endprimitive
// Revision history:
// ----------------
// v1.2  08-Jun-1999  Changing 10ps to 1ps
// v1.1  17-Mar-1999 24 date and time created 99/03/17 17
// v1.2  08-Jun-1999  Changing 10ps to 1ps
// v1.1  17-Mar-1999 24 date and time created 99/03/17 17
// 19 Dec 2006 : Sharavathi : changed the timescale for functiononly option to 
//                            1ns/1ps
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DLY02 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 2.0 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DLY03 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 3.0 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DLY05 (  A , Y );

// Verilog Port Declaration section

   input  A;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           buf #0 TI_BUF_PRIM0 ( Y , A ) ;

`ifdef TI_functiononly
`else

specify

    (A => Y)  = 5.0 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DNC20 (CLK , CLRZ, D, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect


//  Verilog Notifier declaration section

    wire GVCnotifier1 ;
    wire GVCnotifier2 ;

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
           not   TI_NOT_PRIM1 ( IINVnet2, IINVnet1 ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, GVC_D_D, IINVnet2, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, FNET2, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM2 ( IINVnet1, CLK ) ;
           not   TI_NOT_PRIM3 ( IINVnet2, IINVnet1 ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, D, IINVnet2, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( BFONET1, FNET2, IINVnet1, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM4 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM5 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_Q_NOTEQ_D_CLRZ_NOT0_ , Q , GVC_D_D , 1'bx , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif


`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_CLRZ_CLRZ;
    wire TCHKON_AND_Q;
    wire TCHKON_AND_D;
    wire TCHKON_AND_GVC_D_D;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_;
    wire TCHKON_AND_CLRZ;

    and TI_AND_GVC_CLRZ_CLRZ (TCHKON_AND_GVC_CLRZ_CLRZ, GVC_CLRZ_CLRZ, TCHKON_NET);
    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_D (TCHKON_AND_D, D, TCHKON_NET);
    and TI_AND_GVC_D_D (TCHKON_AND_GVC_D_D, GVC_D_D, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_, GVC_Q_NOTEQ_D_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_CLRZ (TCHKON_AND_CLRZ, CLRZ, TCHKON_NET);

`endif


specify

      (CLK  *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK  *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(negedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(negedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge CLRZ,  negedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_D != 0 , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLRZ &&& TCHKON_AND_Q != 0  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.5 11-Sep-2007 :Dundappa.
//                   Added the default delay of 1 for the output pins.
// v1.4 24 Apr 2006 :Sharavathi : Removed TI_veritime options and updated to support 
//                                Simulation without transimiting X when violation
//                                occurs by using Xon
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version
// v2.0 6-oct-2009 Mathangi Updated for non aligned models
// v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DNC40 (CLK , CLRZ, D, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect


//  Verilog Notifier declaration section

    wire GVCnotifier1 ;
    wire GVCnotifier2 ;

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
           not   TI_NOT_PRIM1 ( IINVnet2, IINVnet1 ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, GVC_D_D, IINVnet2, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, FNET2, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM2 ( IINVnet1, CLK ) ;
           not   TI_NOT_PRIM3 ( IINVnet2, IINVnet1 ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, D, IINVnet2, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( BFONET1, FNET2, IINVnet1, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM4 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM5 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_Q_NOTEQ_D_CLRZ_NOT0_ , Q , GVC_D_D , 1'bx , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif


`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_CLRZ_CLRZ;
    wire TCHKON_AND_Q;
    wire TCHKON_AND_D;
    wire TCHKON_AND_GVC_D_D;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_;
    wire TCHKON_AND_CLRZ;

    and TI_AND_GVC_CLRZ_CLRZ (TCHKON_AND_GVC_CLRZ_CLRZ, GVC_CLRZ_CLRZ, TCHKON_NET);
    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_D (TCHKON_AND_D, D, TCHKON_NET);
    and TI_AND_GVC_D_D (TCHKON_AND_GVC_D_D, GVC_D_D, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_, GVC_Q_NOTEQ_D_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_CLRZ (TCHKON_AND_CLRZ, CLRZ, TCHKON_NET);

`endif


specify

      (CLK  *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK  *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(negedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(negedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge CLRZ,  negedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_D != 0 , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLRZ &&& TCHKON_AND_Q != 0  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.5 11-Sep-2007 :Dundappa.
//                   Added the default delay of 1 for the output pins.
// v1.4 24 Apr 2006 :Sharavathi : Removed TI_veritime options and updated to support 
//                                Simulation without transimiting X when violation
//                                occurs by using Xon
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version
// v2.0 6-oct-2009 Mathangi Updated for non aligned models
// v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DTB20 (CLK , CLRZ, D, PREZ, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input PREZ;
   output Q;
   output QZ;
`ifdef TETRAMAX
   _INV I1  ( CLRZ,CLR);
   _INV I2  ( PREZ,PRE);
   _NAND N1 ( CLR,PRE,CLR_PRE);
   _DFF FF1 ( !PREZ, !CLRZ, CLK, D, QINT);
   _INV I3  ( QINT,QZINT);
   _AND A1  ( CLRZ,QINT,Q1);
   _AND A2  ( PRE,CLR_PRE,Q2);
   _AND A3  ( QZINT,PREZ, Q3);
   _AND A4  ( CLR, CLR_PRE, Q4);
   _OR  O1  ( Q1,Q2,Q);
   _OR  O2  ( Q3,Q4,QZ);
`else
`ifdef TI_verilog    
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     parameter Xon = 1;
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);

// Verilog Structure section (in terms of gate prims)

`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ,  GVC_PREZ_PREZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
        dlaudp   TI_DLA_UDP0 ( FNET4, GVC_D_D, IINVnet1, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP1 ( BFONET1, FNET4, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP0 ( BFONET2, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, BFONET1 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
        dlaudp   TI_DLA_UDP2 ( FNET4, D, IINVnet1, CLRZ, PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP3 ( BFONET1, FNET4, CLK, CLRZ, PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP1 ( BFONET2, CLRZ, PREZ, BFONET1 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          buf #1 TI_BUF_PRIM1 ( QZ, BFONET2 ) ;


`else

          buf  TI_BUF_PRIM2 ( Q, BFONET1 ) ;
          buf  TI_BUF_PRIM3 ( QZ, BFONET2 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_CLRZ_NOT0_PREZ_NOT0_ , 1'b0 , 1'b1 , 1'bx , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOT0_PREZ_NOT0_ , 1'b0 , GVC_D_D , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_D_NOT1_CLRZ_NOT0_ , 1'b1 , GVC_D_D , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ , Q , GVC_D_D , 1'bx , 1'b1 , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND4 ( GVC_Q_NOT0_PREZ_NOT0_ , Q , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND5 ( GVC_Q_NOT1_CLRZ_NOT0_ , Q , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif


`ifdef TI_functiononly

specify
    $recovery(posedge PREZ ,posedge CLRZ ,1 , GVCnotifier2_zd );
endspecify

`else
`ifdef TI_verilog

    wire TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_;

    and TI_AND_GVC_D_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_, GVC_D_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_, GVC_Q_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_, GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_, GVC_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_, GVC_D_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_, GVC_Q_NOT1_CLRZ_NOT0_, TCHKON_NET);

`endif


specify
      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

 

`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_ != 0  , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $setuphold(posedge PREZ &&& (TCHKON_NET != 0) , posedge CLRZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_PREZ_PREZ, GVC_CLRZ_CLRZ ); 
   $setuphold(posedge CLRZ &&& (TCHKON_NET != 0) , posedge PREZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ  &&& TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge PREZ  &&& TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

`endif // ifdef TETRAMAX
endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.7 11-Sep-2007 :Dundappa.
//                   Added the default delay of 1 for the output pins.
// v1.6 23-Oct-2002 :Removed `define TI_verilog for 
//                   enabling notiming checks

// v1.5  14-Jan-2002 Modified the timescale 1 ns / 1 ns in TI_functiononly mode to
//                   1 ns/1 ps Track Id 22904
// v1.4  11-Dec-2001 The model is modified by removing conditional paths. For more
//                   information see the Track 23313 TrackId23313
// v1.3  05-Sep-2001 Removed the Copyright block
// v1.2  11-Apr-2000 Updated for Tetramax support
// v1.1  13-Dec-1998 Initial Version
// v2.0  6-oct-2009 Mathangi Updated for non aligned models
// v2.0  9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DTB23 (CLK , CLRZ, D, PREZ, Q ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input PREZ;
   output Q;
`ifdef TETRAMAX
   _INV I1  ( CLRZ,CLR);
   _INV I2  ( PREZ,PRE);
   _NAND N1 ( CLR,PRE,CLR_PRE);
   _DFF FF1 ( !PREZ, !CLRZ, CLK, D, QINT);
   _AND A1  ( CLRZ,QINT,Q1);
   _AND A2  ( PRE,CLR_PRE,Q2);
   _OR  O1  ( Q1,Q2,Q);
`else
`ifdef TI_verilog    
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     parameter Xon = 1;
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);

// Verilog Structure section (in terms of gate prims)

`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ,  GVC_PREZ_PREZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
        dlaudp   TI_DLA_UDP0 ( FNET4, GVC_D_D, IINVnet1, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP1 ( BFONET1, FNET4, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
        dlaudp   TI_DLA_UDP2 ( FNET4, D, IINVnet1, CLRZ, PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP3 ( BFONET1, FNET4, CLK, CLRZ, PREZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;

`else

          buf  TI_BUF_PRIM2 ( Q, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_CLRZ_NOT0_PREZ_NOT0_ , 1'b0 , 1'b1 , 1'bx , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOT0_PREZ_NOT0_ , 1'b0 , GVC_D_D , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_D_NOT1_CLRZ_NOT0_ , 1'b1 , GVC_D_D , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ , Q , GVC_D_D , 1'bx , 1'b1 , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND4 ( GVC_Q_NOT0_PREZ_NOT0_ , Q , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND5 ( GVC_Q_NOT1_CLRZ_NOT0_ , Q , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly

specify
    $recovery(posedge PREZ ,posedge CLRZ ,1 , GVCnotifier2_zd );
endspecify

`else
`ifdef TI_verilog

    wire TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_;

    and TI_AND_GVC_D_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_, GVC_D_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_, GVC_Q_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_, GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_, GVC_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_, GVC_D_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_, GVC_Q_NOT1_CLRZ_NOT0_, TCHKON_NET);

`endif

specify
      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_ != 0  , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $setuphold(posedge PREZ &&& (TCHKON_NET != 0) , posedge CLRZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_PREZ_PREZ, GVC_CLRZ_CLRZ ); 
   $setuphold(posedge CLRZ &&& (TCHKON_NET != 0) , posedge PREZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ  &&& TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge PREZ  &&& TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

`endif // ifdef TETRAMAX
endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------
// v1.7 11-Sep-2007 :Dundappa.
//                   Added the default delay of 1 for the output pins.
// v1.6 23-Oct-2002 :Removed `define TI_verilog for 
//                   enabling notiming checks

// v1.5  14-Jan-2002 Modified the timescale 1 ns / 1 ns in TI_functiononly mode to
//                   1 ns/1 ps Track Id 22904
// v1.4  11-Dec-2001 The model is modified by removing conditional paths. For more
//                   information see the Track 23313 TrackId23313
// v1.3  05-Sep-2001 Removed the Copyright block
// v1.2  11-Apr-2000 Updated for Tetramax support
// v1.1  13-Dec-1998 Initial Version
// v2.0  6-oct-2009  Mathangi Updated for non aligned models
// v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2002 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------


`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DTB24 (CLK , CLRZ, D, PREZ, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input PREZ;
   output QZ;
`ifdef TETRAMAX
   _INV I1  ( CLRZ,CLR);
   _INV I2  ( PREZ,PRE);
   _NAND N1 ( CLR,PRE,CLR_PRE);
   _DFF FF1 ( !PREZ, !CLRZ, CLK, D, QINT);
   _INV I3  ( QINT,QZINT);
   _AND A3  ( QZINT,PREZ, Q3);
   _AND A4  ( CLR, CLR_PRE, Q4);
   _OR  O2  ( Q3,Q4,QZ);
`else
`ifdef TI_verilog    
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     parameter Xon = 1;
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ,  GVC_PREZ_PREZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
        dlaudp   TI_DLA_UDP0 ( FNET4, GVC_D_D, IINVnet1, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP1 ( BFONET1, FNET4, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP0 ( BFONET2, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, BFONET1 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
        dlaudp   TI_DLA_UDP2 ( FNET4, D, IINVnet1, CLRZ, PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP3 ( BFONET1, FNET4, CLK, CLRZ, PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP1 ( BFONET2, CLRZ, PREZ, BFONET1 ) ;


`endif

`ifdef TI_functiononly

           not    TI_BUF_PRIM0 ( NOT_QZ, QZ ) ;
           buf #1 TI_BUF_PRIM1 ( QZ, BFONET2 ) ;

`else
           not   TI_BUF_PRIM1 ( NOT_QZ, QZ ) ;
           buf  TI_BUF_PRIM3 ( QZ, BFONET2 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_CLRZ_NOT0_PREZ_NOT0_ , 1'b0 , 1'b1 , 1'bx , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOT0_PREZ_NOT0_ , 1'b0 , GVC_D_D , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_D_NOT1_CLRZ_NOT0_ , 1'b1 , GVC_D_D , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ , NOT_QZ , GVC_D_D , 1'bx , 1'b1 , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND4 ( GVC_Q_NOT0_PREZ_NOT0_ , NOT_QZ , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND5 ( GVC_Q_NOT1_CLRZ_NOT0_ , NOT_QZ , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif


`ifdef TI_functiononly

specify
    $recovery(posedge PREZ ,posedge CLRZ ,1 , GVCnotifier2_zd );
endspecify

`else
`ifdef TI_verilog

    wire TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_;

    and TI_AND_GVC_D_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_, GVC_D_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_, GVC_Q_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_, GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_, GVC_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_, GVC_D_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_, GVC_Q_NOT1_CLRZ_NOT0_, TCHKON_NET);

`endif


specify
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ != 0 ) , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ != 0 ) , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_ != 0 ) , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_ != 0 ) , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $setuphold(posedge PREZ &&& (TCHKON_NET != 0) , posedge CLRZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_PREZ_PREZ, GVC_CLRZ_CLRZ ); 
   $setuphold(posedge CLRZ &&& (TCHKON_NET != 0) , posedge PREZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ ); 
   $width(posedge CLK  &&& ( TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ != 0 )  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& ( TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ != 0 )  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ  &&& ( TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_ != 0 )  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge PREZ  &&& ( TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_ != 0 )  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

`endif // ifdef TETRAMAX
endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.7 11-Sep-2007 :Dundappa.
//                   Added the default delay of 1 for the output pins.
// v1.6 23-Oct-2002 :Removed `define TI_verilog for 
//                   enabling notiming checks

// v1.5  14-Jan-2002 Modified the timescale 1 ns / 1 ns in TI_functiononly mode to
//                   1 ns/1 ps Track Id 22904
// v1.4  11-Dec-2001 The model is modified by removing conditional paths. For more
//                   information see the Track 23313 TrackId23313
// v1.3  05-Sep-2001 Removed the Copyright block
// v1.2  11-Apr-2000 Updated for Tetramax support
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//    22-Jan-2010 Mazhar. Added TCHKON_NET switch for setuphold
//                of prez <---> clrz paths
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DTB40 (CLK , CLRZ, D, PREZ, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input PREZ;
   output Q;
   output QZ;
`ifdef TETRAMAX
   _INV I1  ( CLRZ,CLR);
   _INV I2  ( PREZ,PRE);
   _NAND N1 ( CLR,PRE,CLR_PRE);
   _DFF FF1 ( !PREZ, !CLRZ, CLK, D, QINT);
   _INV I3  ( QINT,QZINT);
   _AND A1  ( CLRZ,QINT,Q1);
   _AND A2  ( PRE,CLR_PRE,Q2);
   _AND A3  ( QZINT,PREZ, Q3);
   _AND A4  ( CLR, CLR_PRE, Q4);
   _OR  O1  ( Q1,Q2,Q);
   _OR  O2  ( Q3,Q4,QZ);
`else
`ifdef TI_verilog    
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     parameter Xon = 1;
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);

// Verilog Structure section (in terms of gate prims)

`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ,  GVC_PREZ_PREZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
        dlaudp   TI_DLA_UDP0 ( FNET4, GVC_D_D, IINVnet1, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP1 ( BFONET1, FNET4, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP0 ( BFONET2, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, BFONET1 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
        dlaudp   TI_DLA_UDP2 ( FNET4, D, IINVnet1, CLRZ, PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP3 ( BFONET1, FNET4, CLK, CLRZ, PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP1 ( BFONET2, CLRZ, PREZ, BFONET1 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          buf #1 TI_BUF_PRIM1 ( QZ, BFONET2 ) ;


`else

          buf  TI_BUF_PRIM2 ( Q, BFONET1 ) ;
          buf  TI_BUF_PRIM3 ( QZ, BFONET2 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_CLRZ_NOT0_PREZ_NOT0_ , 1'b0 , 1'b1 , 1'bx , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOT0_PREZ_NOT0_ , 1'b0 , GVC_D_D , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_D_NOT1_CLRZ_NOT0_ , 1'b1 , GVC_D_D , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ , Q , GVC_D_D , 1'bx , 1'b1 , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND4 ( GVC_Q_NOT0_PREZ_NOT0_ , Q , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND5 ( GVC_Q_NOT1_CLRZ_NOT0_ , Q , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif


`ifdef TI_functiononly

specify
    $recovery(posedge PREZ ,posedge CLRZ ,1 , GVCnotifier2_zd );
endspecify

`else
`ifdef TI_verilog

    wire TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_;

    and TI_AND_GVC_D_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_, GVC_D_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_, GVC_Q_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_, GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_, GVC_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_, GVC_D_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_, GVC_Q_NOT1_CLRZ_NOT0_, TCHKON_NET);

`endif


specify
      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

 

`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_ != 0  , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $setuphold(posedge PREZ &&& (TCHKON_NET != 0) , posedge CLRZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_PREZ_PREZ, GVC_CLRZ_CLRZ ); 
   $setuphold(posedge CLRZ &&& (TCHKON_NET != 0) , posedge PREZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ  &&& TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge PREZ  &&& TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

`endif // ifdef TETRAMAX
endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.7 11-Sep-2007 :Dundappa.
//                   Added the default delay of 1 for the output pins.
// v1.6 23-Oct-2002 :Removed `define TI_verilog for 
//                   enabling notiming checks

// v1.5  14-Jan-2002 Modified the timescale 1 ns / 1 ns in TI_functiononly mode to
//                   1 ns/1 ps Track Id 22904
// v1.4  11-Dec-2001 The model is modified by removing conditional paths. For more
//                   information see the Track 23313 TrackId23313
// v1.3  05-Sep-2001 Removed the Copyright block
// v1.2  11-Apr-2000 Updated for Tetramax support
// v1.1  13-Dec-1998 Initial Version
// v2.0  6-oct-2009 Mathangi Updated for non aligned models
// v2.0  9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DTB43 (CLK , CLRZ, D, PREZ, Q ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input PREZ;
   output Q;
`ifdef TETRAMAX
   _INV I1  ( CLRZ,CLR);
   _INV I2  ( PREZ,PRE);
   _NAND N1 ( CLR,PRE,CLR_PRE);
   _DFF FF1 ( !PREZ, !CLRZ, CLK, D, QINT);
   _AND A1  ( CLRZ,QINT,Q1);
   _AND A2  ( PRE,CLR_PRE,Q2);
   _OR  O1  ( Q1,Q2,Q);
`else
`ifdef TI_verilog    
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     parameter Xon = 1;
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);

// Verilog Structure section (in terms of gate prims)

`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ,  GVC_PREZ_PREZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
        dlaudp   TI_DLA_UDP0 ( FNET4, GVC_D_D, IINVnet1, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP1 ( BFONET1, FNET4, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
        dlaudp   TI_DLA_UDP2 ( FNET4, D, IINVnet1, CLRZ, PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP3 ( BFONET1, FNET4, CLK, CLRZ, PREZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;

`else

          buf  TI_BUF_PRIM2 ( Q, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_CLRZ_NOT0_PREZ_NOT0_ , 1'b0 , 1'b1 , 1'bx , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOT0_PREZ_NOT0_ , 1'b0 , GVC_D_D , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_D_NOT1_CLRZ_NOT0_ , 1'b1 , GVC_D_D , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ , Q , GVC_D_D , 1'bx , 1'b1 , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND4 ( GVC_Q_NOT0_PREZ_NOT0_ , Q , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND5 ( GVC_Q_NOT1_CLRZ_NOT0_ , Q , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly

specify
    $recovery(posedge PREZ ,posedge CLRZ ,1 , GVCnotifier2_zd );
endspecify

`else
`ifdef TI_verilog

    wire TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_;

    and TI_AND_GVC_D_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_, GVC_D_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_, GVC_Q_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_, GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_, GVC_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_, GVC_D_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_, GVC_Q_NOT1_CLRZ_NOT0_, TCHKON_NET);

`endif

specify
      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_ != 0  , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $setuphold(posedge PREZ &&& (TCHKON_NET != 0) , posedge CLRZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_PREZ_PREZ, GVC_CLRZ_CLRZ ); 
   $setuphold(posedge CLRZ &&& (TCHKON_NET != 0) , posedge PREZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ  &&& TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge PREZ  &&& TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

`endif // ifdef TETRAMAX
endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------
// v1.7 11-Sep-2007 :Dundappa.
//                   Added the default delay of 1 for the output pins.
// v1.6 23-Oct-2002 :Removed `define TI_verilog for 
//                   enabling notiming checks

// v1.5  14-Jan-2002 Modified the timescale 1 ns / 1 ns in TI_functiononly mode to
//                   1 ns/1 ps Track Id 22904
// v1.4  11-Dec-2001 The model is modified by removing conditional paths. For more
//                   information see the Track 23313 TrackId23313
// v1.3  05-Sep-2001 Removed the Copyright block
// v1.2  11-Apr-2000 Updated for Tetramax support
// v1.1  13-Dec-1998 Initial Version
// v2.0  6-oct-2009  Mathangi Updated for non aligned models
// v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2002 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------


`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DTB44 (CLK , CLRZ, D, PREZ, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input PREZ;
   output QZ;
`ifdef TETRAMAX
   _INV I1  ( CLRZ,CLR);
   _INV I2  ( PREZ,PRE);
   _NAND N1 ( CLR,PRE,CLR_PRE);
   _DFF FF1 ( !PREZ, !CLRZ, CLK, D, QINT);
   _INV I3  ( QINT,QZINT);
   _AND A3  ( QZINT,PREZ, Q3);
   _AND A4  ( CLR, CLR_PRE, Q4);
   _OR  O2  ( Q3,Q4,QZ);
`else
`ifdef TI_verilog    
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     parameter Xon = 1;
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ,  GVC_PREZ_PREZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
        dlaudp   TI_DLA_UDP0 ( FNET4, GVC_D_D, IINVnet1, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP1 ( BFONET1, FNET4, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP0 ( BFONET2, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, BFONET1 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
        dlaudp   TI_DLA_UDP2 ( FNET4, D, IINVnet1, CLRZ, PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP3 ( BFONET1, FNET4, CLK, CLRZ, PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP1 ( BFONET2, CLRZ, PREZ, BFONET1 ) ;


`endif

`ifdef TI_functiononly

           not    TI_BUF_PRIM0 ( NOT_QZ, QZ ) ;
           buf #1 TI_BUF_PRIM1 ( QZ, BFONET2 ) ;

`else
           not   TI_BUF_PRIM1 ( NOT_QZ, QZ ) ;
           buf  TI_BUF_PRIM3 ( QZ, BFONET2 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_CLRZ_NOT0_PREZ_NOT0_ , 1'b0 , 1'b1 , 1'bx , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOT0_PREZ_NOT0_ , 1'b0 , GVC_D_D , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_D_NOT1_CLRZ_NOT0_ , 1'b1 , GVC_D_D , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ , NOT_QZ , GVC_D_D , 1'bx , 1'b1 , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND4 ( GVC_Q_NOT0_PREZ_NOT0_ , NOT_QZ , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND5 ( GVC_Q_NOT1_CLRZ_NOT0_ , NOT_QZ , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif


`ifdef TI_functiononly

specify
    $recovery(posedge PREZ ,posedge CLRZ ,1 , GVCnotifier2_zd );
endspecify

`else
`ifdef TI_verilog

    wire TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_;

    and TI_AND_GVC_D_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_, GVC_D_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_, GVC_Q_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_, GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_, GVC_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_, GVC_D_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_, GVC_Q_NOT1_CLRZ_NOT0_, TCHKON_NET);

`endif


specify
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ != 0 ) , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ != 0 ) , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_ != 0 ) , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_ != 0 ) , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $setuphold(posedge PREZ &&& (TCHKON_NET != 0) , posedge CLRZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_PREZ_PREZ, GVC_CLRZ_CLRZ ); 
   $setuphold(posedge CLRZ &&& (TCHKON_NET != 0) , posedge PREZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ ); 
   $width(posedge CLK  &&& ( TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ != 0 )  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& ( TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_PREZ_NOT0_ != 0 )  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ  &&& ( TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_ != 0 )  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge PREZ  &&& ( TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_ != 0 )  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

`endif // ifdef TETRAMAX
endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.7 11-Sep-2007 :Dundappa.
//                   Added the default delay of 1 for the output pins.
// v1.6 23-Oct-2002 :Removed `define TI_verilog for 
//                   enabling notiming checks

// v1.5  14-Jan-2002 Modified the timescale 1 ns / 1 ns in TI_functiononly mode to
//                   1 ns/1 ps Track Id 22904
// v1.4  11-Dec-2001 The model is modified by removing conditional paths. For more
//                   information see the Track 23313 TrackId23313
// v1.3  05-Sep-2001 Removed the Copyright block
// v1.2  11-Apr-2000 Updated for Tetramax support
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//    22-Jan-2010 Mazhar. Added TCHKON_NET switch for setuphold
//                of prez <---> clrz paths
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DTC20 (CLK , CLRZ, D, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   output Q;
   output QZ;

`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, D, IINVnet1, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( BFONET1, FNET2, CLK, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_Q_NOTEQ_D_CLRZ_NOT0_ , Q , GVC_D_D , 1'bx , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else
`ifdef TI_verilog

    wire TCHKON_AND_GVC_CLRZ_CLRZ;
    wire TCHKON_AND_Q;
    wire TCHKON_AND_D;
    wire TCHKON_AND_GVC_D_D;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_;
    wire TCHKON_AND_CLRZ;

    and TI_AND_GVC_CLRZ_CLRZ (TCHKON_AND_GVC_CLRZ_CLRZ, GVC_CLRZ_CLRZ, TCHKON_NET);
    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_D (TCHKON_AND_D, D, TCHKON_NET);
    and TI_AND_GVC_D_D (TCHKON_AND_GVC_D_D, GVC_D_D, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_, GVC_Q_NOTEQ_D_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_CLRZ (TCHKON_AND_CLRZ, CLRZ, TCHKON_NET);

`endif


specify

      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_D != 0 , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& TCHKON_AND_Q != 0  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.6 11-Sep-2007 :Dundappa.
//                   Added the default delay of 1 for the output pins.
// v1.5 23-Oct-2002 :Removed `define TI_verilog for 
//                   enabling notiming checks

// v1.4  14-Jan-2002 Modified the timescale 1 ns / 1 ns in TI_functiononly mode to
//                   1 ns/1 ps Track Id 22904
// v1.3  11-Dec-2001 The model is modified by removing conditional paths. For more
//                   information see the Track 23313 TrackId23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module DTC21 (CLK , CLRZ, D, LD, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input LD;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ,  GVC_LD_LD  ; 

           not   TI_NOT_PRIM0 (NOT_GVC_LD_LD , GVC_LD_LD ) ;
        mu1udp   TI_MUX2_UDP0 ( DIN, NOT_GVC_LD_LD, GVC_D_D, BFONET1 ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, GVC_CLK_CLK ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, DIN, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM2 ( NOT_LD, LD ) ;
        mu1udp   TI_MUX2_UDP1 ( DIN, NOT_LD, D, BFONET1 ) ;
           not   TI_NOT_PRIM3 ( IINVnet1, CLK ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, DIN, IINVnet1, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( BFONET1, FNET2, CLK, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM4 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM5 ( QZ, BFONET1 ) ;
 
 
`else
 
          buf  TI_BUF_PRIM6 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM7 ( QZ, BFONET1 ) ;



`endif
 
`ifdef TI_verilog
 
//  Logic enabling constraint check statements for verilog/verifault
 
      //  not TI_NOT_PRIM4 ( NOT_ENZ, GVC_ENZ_ENZ ) ;
        and TI_AND_PRIM0 ( GVC_LD_NOT0_CLRZ_NOT0_ , GVC_LD_LD , GVC_CLRZ_CLRZ ) ;
        xor TI_XOR_PRIM0 ( D_NOTEQ_Q , GVC_D_D , Q ) ;
        and TI_AND_PRIM1 ( GVC_D_NOTEQ_Q_CLRZ_NOT0_ , D_NOTEQ_Q , GVC_CLRZ_CLRZ ) ;
        and TI_AND_PRIM2 ( GVC_D_NOT0_LD_NOT0_, GVC_D_D, GVC_LD_LD ) ;
        and TI_AND_PRIM3 ( GVC_Q_NOTEQ_D_CLRZ_NOT0_LD_NOT0_ , D_NOTEQ_Q , GVC_CLRZ_CLRZ , GVC_LD_LD ) ;
 
`endif
       
 

`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_Q;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_LD_NOT0_;
    wire TCHKON_AND_GVC_D_NOT0_LD_NOT0_;
    wire TCHKON_AND_GVC_LD_NOT0_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0_;

    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_LD_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_LD_NOT0_, GVC_Q_NOTEQ_D_CLRZ_NOT0_LD_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOT0_LD_NOT0_ (TCHKON_AND_GVC_D_NOT0_LD_NOT0_, GVC_D_NOT0_LD_NOT0_, TCHKON_NET);
    and TI_AND_GVC_LD_NOT0_CLRZ_NOT0_ (TCHKON_AND_GVC_LD_NOT0_CLRZ_NOT0_, GVC_LD_NOT0_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0_, GVC_D_NOTEQ_Q_CLRZ_NOT0_, TCHKON_NET);

`endif


specify

      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, TCHKON_AND_GVC_LD_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, TCHKON_AND_GVC_LD_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, TCHKON_AND_GVC_D_NOT0_LD_NOT0_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $setuphold(posedge CLK,  posedge LD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, TCHKON_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_LD_LD ); 
   $setuphold(posedge CLK,  negedge LD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, TCHKON_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_LD_LD ); 
   $width(posedge CLK &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_LD_NOT0_ != 0   ,0.01 : 0.01 : 0.01 ,  0 , GVCnotifier2_zd) ; 
   $width(negedge CLK &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_LD_NOT0_ != 0   ,0.01 : 0.01 : 0.01 ,  0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& TCHKON_AND_Q != 0   ,0.01 : 0.01 : 0.01 ,  0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.3 11-Sep-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.2  18-Sep-1999 Duplicate instance names were corrected
// v1.1  03-Sep-1999 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DTC23 (CLK , CLRZ, D, Q ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   output Q;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, D, IINVnet1, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( BFONET1, FNET2, CLK, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_Q_NOTEQ_D_CLRZ_NOT0_ , Q , GVC_D_D , 1'bx , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif


`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_CLRZ_CLRZ;
    wire TCHKON_AND_Q;
    wire TCHKON_AND_D;
    wire TCHKON_AND_GVC_D_D;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_;
    wire TCHKON_AND_CLRZ;

    and TI_AND_GVC_CLRZ_CLRZ (TCHKON_AND_GVC_CLRZ_CLRZ, GVC_CLRZ_CLRZ, TCHKON_NET);
    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_D (TCHKON_AND_D, D, TCHKON_NET);
    and TI_AND_GVC_D_D (TCHKON_AND_GVC_D_D, GVC_D_D, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_, GVC_Q_NOTEQ_D_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_CLRZ (TCHKON_AND_CLRZ, CLRZ, TCHKON_NET);

`endif


specify

      (CLK  *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_D != 0 , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& TCHKON_AND_Q != 0  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module DTC24 (CLK , CLRZ, D, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( Q, FNET2, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, D, IINVnet1, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( Q, FNET2, CLK, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          not #1 TI_NOT_PRIM2 ( QZ, Q ) ;


`else

          not  TI_NOT_PRIM3 ( QZ, Q ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    not TI_NOT_PRIM4 (GVCnet0 , GVC_D_D);
    cons_udp TI_COND0 ( GVC_QZ_NOTEQ_D_CLRZ_NOT0_ , QZ , GVCnet0 , 1'bx , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_CLRZ_CLRZ;
    wire TCHKON_AND_GVC_QZ_NOTEQ_D_CLRZ_NOT0_;
    wire TCHKON_AND_D;
    wire TCHKON_AND_GVC_D_D;
    wire TCHKON_AND_CLRZ;

    and TI_AND_GVC_CLRZ_CLRZ (TCHKON_AND_GVC_CLRZ_CLRZ, GVC_CLRZ_CLRZ, TCHKON_NET);
    and TI_AND_GVC_QZ_NOTEQ_D_CLRZ_NOT0_ (TCHKON_AND_GVC_QZ_NOTEQ_D_CLRZ_NOT0_, GVC_QZ_NOTEQ_D_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_D (TCHKON_AND_D, D, TCHKON_NET);
    and TI_AND_GVC_D_D (TCHKON_AND_GVC_D_D, GVC_D_D, TCHKON_NET);
    and TI_AND_CLRZ (TCHKON_AND_CLRZ, CLRZ, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_QZ;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_QZ (NOT_TCHKON_OR_QZ, QZ, TCHKON_INV);

`endif


specify

      (CLK  *> QZ  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);



`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_D != 0 , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& NOT_TCHKON_OR_QZ != 1  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DTC40 (CLK , CLRZ, D, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   output Q;
   output QZ;

`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, D, IINVnet1, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( BFONET1, FNET2, CLK, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_Q_NOTEQ_D_CLRZ_NOT0_ , Q , GVC_D_D , 1'bx , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else
`ifdef TI_verilog

    wire TCHKON_AND_GVC_CLRZ_CLRZ;
    wire TCHKON_AND_Q;
    wire TCHKON_AND_D;
    wire TCHKON_AND_GVC_D_D;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_;
    wire TCHKON_AND_CLRZ;

    and TI_AND_GVC_CLRZ_CLRZ (TCHKON_AND_GVC_CLRZ_CLRZ, GVC_CLRZ_CLRZ, TCHKON_NET);
    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_D (TCHKON_AND_D, D, TCHKON_NET);
    and TI_AND_GVC_D_D (TCHKON_AND_GVC_D_D, GVC_D_D, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_, GVC_Q_NOTEQ_D_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_CLRZ (TCHKON_AND_CLRZ, CLRZ, TCHKON_NET);

`endif


specify

      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_D != 0 , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& TCHKON_AND_Q != 0  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.6 11-Sep-2007 :Dundappa.
//                   Added the default delay of 1 for the output pins.
// v1.5 23-Oct-2002 :Removed `define TI_verilog for 
//                   enabling notiming checks

// v1.4  14-Jan-2002 Modified the timescale 1 ns / 1 ns in TI_functiononly mode to
//                   1 ns/1 ps Track Id 22904
// v1.3  11-Dec-2001 The model is modified by removing conditional paths. For more
//                   information see the Track 23313 TrackId23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module DTC41 (CLK , CLRZ, D, LD, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input LD;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ,  GVC_LD_LD  ; 

           not   TI_NOT_PRIM0 (NOT_GVC_LD_LD , GVC_LD_LD ) ;
        mu1udp   TI_MUX2_UDP0 ( DIN, NOT_GVC_LD_LD, GVC_D_D, BFONET1 ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, GVC_CLK_CLK ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, DIN, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM2 ( NOT_LD, LD ) ;
        mu1udp   TI_MUX2_UDP1 ( DIN, NOT_LD, D, BFONET1 ) ;
           not   TI_NOT_PRIM3 ( IINVnet1, CLK ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, DIN, IINVnet1, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( BFONET1, FNET2, CLK, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM4 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM5 ( QZ, BFONET1 ) ;
 
 
`else
 
          buf  TI_BUF_PRIM6 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM7 ( QZ, BFONET1 ) ;



`endif
 
`ifdef TI_verilog
 
//  Logic enabling constraint check statements for verilog/verifault
 
      //  not TI_NOT_PRIM4 ( NOT_ENZ, GVC_ENZ_ENZ ) ;
        and TI_AND_PRIM0 ( GVC_LD_NOT0_CLRZ_NOT0_ , GVC_LD_LD , GVC_CLRZ_CLRZ ) ;
        xor TI_XOR_PRIM0 ( D_NOTEQ_Q , GVC_D_D , Q ) ;
        and TI_AND_PRIM1 ( GVC_D_NOTEQ_Q_CLRZ_NOT0_ , D_NOTEQ_Q , GVC_CLRZ_CLRZ ) ;
        and TI_AND_PRIM2 ( GVC_D_NOT0_LD_NOT0_, GVC_D_D, GVC_LD_LD ) ;
        and TI_AND_PRIM3 ( GVC_Q_NOTEQ_D_CLRZ_NOT0_LD_NOT0_ , D_NOTEQ_Q , GVC_CLRZ_CLRZ , GVC_LD_LD ) ;
 
`endif
       
 

`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_Q;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_LD_NOT0_;
    wire TCHKON_AND_GVC_D_NOT0_LD_NOT0_;
    wire TCHKON_AND_GVC_LD_NOT0_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0_;

    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_LD_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_LD_NOT0_, GVC_Q_NOTEQ_D_CLRZ_NOT0_LD_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOT0_LD_NOT0_ (TCHKON_AND_GVC_D_NOT0_LD_NOT0_, GVC_D_NOT0_LD_NOT0_, TCHKON_NET);
    and TI_AND_GVC_LD_NOT0_CLRZ_NOT0_ (TCHKON_AND_GVC_LD_NOT0_CLRZ_NOT0_, GVC_LD_NOT0_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0_, GVC_D_NOTEQ_Q_CLRZ_NOT0_, TCHKON_NET);

`endif


specify

      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, TCHKON_AND_GVC_LD_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, TCHKON_AND_GVC_LD_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, TCHKON_AND_GVC_D_NOT0_LD_NOT0_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $setuphold(posedge CLK,  posedge LD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, TCHKON_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_LD_LD ); 
   $setuphold(posedge CLK,  negedge LD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, TCHKON_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_LD_LD ); 
   $width(posedge CLK &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_LD_NOT0_ != 0   ,0.01 : 0.01 : 0.01 ,  0 , GVCnotifier2_zd) ; 
   $width(negedge CLK &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_LD_NOT0_ != 0   ,0.01 : 0.01 : 0.01 ,  0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& TCHKON_AND_Q != 0   ,0.01 : 0.01 : 0.01 ,  0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.3 11-Sep-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.2  18-Sep-1999 Duplicate instance names were corrected
// v1.1  03-Sep-1999 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DTC43 (CLK , CLRZ, D, Q ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   output Q;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, D, IINVnet1, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( BFONET1, FNET2, CLK, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_Q_NOTEQ_D_CLRZ_NOT0_ , Q , GVC_D_D , 1'bx , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif


`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_CLRZ_CLRZ;
    wire TCHKON_AND_Q;
    wire TCHKON_AND_D;
    wire TCHKON_AND_GVC_D_D;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_;
    wire TCHKON_AND_CLRZ;

    and TI_AND_GVC_CLRZ_CLRZ (TCHKON_AND_GVC_CLRZ_CLRZ, GVC_CLRZ_CLRZ, TCHKON_NET);
    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_D (TCHKON_AND_D, D, TCHKON_NET);
    and TI_AND_GVC_D_D (TCHKON_AND_GVC_D_D, GVC_D_D, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_, GVC_Q_NOTEQ_D_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_CLRZ (TCHKON_AND_CLRZ, CLRZ, TCHKON_NET);

`endif


specify

      (CLK  *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_D != 0 , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& TCHKON_AND_Q != 0  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module DTC44 (CLK , CLRZ, D, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( Q, FNET2, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, D, IINVnet1, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( Q, FNET2, CLK, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          not #1 TI_NOT_PRIM2 ( QZ, Q ) ;


`else

          not  TI_NOT_PRIM3 ( QZ, Q ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    not TI_NOT_PRIM4 (GVCnet0 , GVC_D_D);
    cons_udp TI_COND0 ( GVC_QZ_NOTEQ_D_CLRZ_NOT0_ , QZ , GVCnet0 , 1'bx , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_CLRZ_CLRZ;
    wire TCHKON_AND_GVC_QZ_NOTEQ_D_CLRZ_NOT0_;
    wire TCHKON_AND_D;
    wire TCHKON_AND_GVC_D_D;
    wire TCHKON_AND_CLRZ;

    and TI_AND_GVC_CLRZ_CLRZ (TCHKON_AND_GVC_CLRZ_CLRZ, GVC_CLRZ_CLRZ, TCHKON_NET);
    and TI_AND_GVC_QZ_NOTEQ_D_CLRZ_NOT0_ (TCHKON_AND_GVC_QZ_NOTEQ_D_CLRZ_NOT0_, GVC_QZ_NOTEQ_D_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_D (TCHKON_AND_D, D, TCHKON_NET);
    and TI_AND_GVC_D_D (TCHKON_AND_GVC_D_D, GVC_D_D, TCHKON_NET);
    and TI_AND_CLRZ (TCHKON_AND_CLRZ, CLRZ, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_QZ;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_QZ (NOT_TCHKON_OR_QZ, QZ, TCHKON_INV);

`endif


specify

      (CLK  *> QZ  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);



`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_D != 0 , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& NOT_TCHKON_OR_QZ != 1  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DTN20 (CLK , D, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_nudp   TI_LACTHN_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_nudp   TI_LACTHN_UDP2 ( FNET2, D, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP3 ( BFONET1, FNET2, CLK, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_Q_NOTEQ_D_ , Q , GVC_D_D , 1'bx , 1'b1 , 1'b1 , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_Q_NOTEQ_D_;

    and TI_AND_GVC_Q_NOTEQ_D_ (TCHKON_AND_GVC_Q_NOTEQ_D_, GVC_Q_NOTEQ_D_, TCHKON_NET);

`endif


specify
    
      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK &&& (TCHKON_NET != 0) ,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK &&& (TCHKON_NET != 0) ,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_D_D ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.5 11-Sep-2007 :Dundappa.
//                   Added the default delay of 1 for the output pins.

// v1.4 23-Oct-2002 :Removed `define TI_verilog for 
//                   enabling notiming checks

// v1.3  14-Jan-2002 Modified the timescale 1 ns / 1 ns in TI_functiononly mode to
//                   1 ns/1 ps Track Id 22904
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models
//v2.0 9-oct-2009 Mathangi Changed 
//     (posedge CLK *> (Q  +: D)) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
//     (posedge CLK *> (QZ  -: D)) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
//to
//    (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
//    (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
// in consistence with the asic model.
  


//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DTN21 (CLK , D, Q ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   output Q;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_nudp   TI_LACTHN_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_nudp   TI_LACTHN_UDP2 ( FNET2, D, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP3 ( BFONET1, FNET2, CLK, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_Q_NOTEQ_D_ , Q , GVC_D_D , 1'bx , 1'b1 , 1'b1 , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_Q_NOTEQ_D_;

    and TI_AND_GVC_Q_NOTEQ_D_ (TCHKON_AND_GVC_Q_NOTEQ_D_, GVC_Q_NOTEQ_D_, TCHKON_NET);

`endif


specify

     (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK &&& (TCHKON_NET != 0) ,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK &&& (TCHKON_NET != 0) ,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_D_D ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.3 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models
//v2.0 9-oct-2009 Mathangi Changed 
//    (posedge CLK *> (Q  +: D)) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
//    to
//    (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
//    in consistence with the asic model.
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DTN22 (CLK , D, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_nudp   TI_LACTHN_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP1 ( Q, FNET2, GVC_CLK_CLK, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_nudp   TI_LACTHN_UDP2 ( FNET2, D, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP3 ( Q, FNET2, CLK, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          not #1 TI_NOT_PRIM2 ( QZ, Q ) ;


`else

          not  TI_NOT_PRIM3 ( QZ, Q ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    not TI_NOT_PRIM4 (GVCnet0 , GVC_D_D);
    cons_udp TI_COND0 ( GVC_QZ_NOTEQ_D_ , QZ , GVCnet0 , 1'bx , 1'b1 , 1'b1 , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_QZ_NOTEQ_D_;

    and TI_AND_GVC_QZ_NOTEQ_D_ (TCHKON_AND_GVC_QZ_NOTEQ_D_, GVC_QZ_NOTEQ_D_, TCHKON_NET);

`endif


specify

     
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK &&& (TCHKON_NET != 0) ,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK &&& (TCHKON_NET != 0) ,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_D_D ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.3 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models
//v2.0 9-oct-2009 Mathangi Changed
//(posedge CLK *> (QZ  -: D)) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
//to
//(CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
// in consistence with the asic model.
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DTN40 (CLK , D, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_nudp   TI_LACTHN_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_nudp   TI_LACTHN_UDP2 ( FNET2, D, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP3 ( BFONET1, FNET2, CLK, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_Q_NOTEQ_D_ , Q , GVC_D_D , 1'bx , 1'b1 , 1'b1 , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_Q_NOTEQ_D_;

    and TI_AND_GVC_Q_NOTEQ_D_ (TCHKON_AND_GVC_Q_NOTEQ_D_, GVC_Q_NOTEQ_D_, TCHKON_NET);

`endif


specify
    
      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK &&& (TCHKON_NET != 0) ,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK &&& (TCHKON_NET != 0) ,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_D_D ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.5 11-Sep-2007 :Dundappa.
//                   Added the default delay of 1 for the output pins.

// v1.4 23-Oct-2002 :Removed `define TI_verilog for 
//                   enabling notiming checks

// v1.3  14-Jan-2002 Modified the timescale 1 ns / 1 ns in TI_functiononly mode to
//                   1 ns/1 ps Track Id 22904
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models
//v2.0 9-oct-2009 Mathangi Changed 
//     (posedge CLK *> (Q  +: D)) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
//     (posedge CLK *> (QZ  -: D)) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
//to
//    (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
//    (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
// in consistence with the asic model.
  


//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DTN41 (CLK , D, Q ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   output Q;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_nudp   TI_LACTHN_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_nudp   TI_LACTHN_UDP2 ( FNET2, D, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP3 ( BFONET1, FNET2, CLK, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_Q_NOTEQ_D_ , Q , GVC_D_D , 1'bx , 1'b1 , 1'b1 , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_Q_NOTEQ_D_;

    and TI_AND_GVC_Q_NOTEQ_D_ (TCHKON_AND_GVC_Q_NOTEQ_D_, GVC_Q_NOTEQ_D_, TCHKON_NET);

`endif


specify

     (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK &&& (TCHKON_NET != 0) ,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK &&& (TCHKON_NET != 0) ,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_D_D ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.3 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models
//v2.0 9-oct-2009 Mathangi Changed 
//    (posedge CLK *> (Q  +: D)) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
//    to
//    (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
//    in consistence with the asic model.
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module DTN42 (CLK , D, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_nudp   TI_LACTHN_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP1 ( Q, FNET2, GVC_CLK_CLK, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_nudp   TI_LACTHN_UDP2 ( FNET2, D, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP3 ( Q, FNET2, CLK, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          not #1 TI_NOT_PRIM2 ( QZ, Q ) ;


`else

          not  TI_NOT_PRIM3 ( QZ, Q ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    not TI_NOT_PRIM4 (GVCnet0 , GVC_D_D);
    cons_udp TI_COND0 ( GVC_QZ_NOTEQ_D_ , QZ , GVCnet0 , 1'bx , 1'b1 , 1'b1 , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_QZ_NOTEQ_D_;

    and TI_AND_GVC_QZ_NOTEQ_D_ (TCHKON_AND_GVC_QZ_NOTEQ_D_, GVC_QZ_NOTEQ_D_, TCHKON_NET);

`endif


specify

     
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK &&& (TCHKON_NET != 0) ,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK &&& (TCHKON_NET != 0) ,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_CLK_CLK, GVC_D_D ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.3 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models
//v2.0 9-oct-2009 Mathangi Changed
//(posedge CLK *> (QZ  -: D)) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
//to
//(CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
// in consistence with the asic model.
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module DTP20 (CLK , D, PREZ, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input PREZ;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_PREZ_PREZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_pudp   TI_LACTHP_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVC_PREZ_PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_PREZ_PREZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_pudp   TI_LACTHP_UDP2 ( FNET2, D, IINVnet1, PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP3 ( BFONET1, FNET2, CLK, PREZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_Q_NOTEQ_D_PREZ_NOT0_ , Q , GVC_D_D , 1'bx , 1'b1 , 1'b1 , GVC_PREZ_PREZ ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_PREZ;
    wire TCHKON_AND_GVC_PREZ_PREZ;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_;

    and TI_AND_PREZ (TCHKON_AND_PREZ, PREZ, TCHKON_NET);
    and TI_AND_GVC_PREZ_PREZ (TCHKON_AND_GVC_PREZ_PREZ, GVC_PREZ_PREZ, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_, GVC_Q_NOTEQ_D_PREZ_NOT0_, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_Q;
    wire NOT_TCHKON_OR_D;
    wire NOT_TCHKON_OR_GVC_D_D;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_Q (NOT_TCHKON_OR_Q, Q, TCHKON_INV);
    or TI_OR_D (NOT_TCHKON_OR_D, D, TCHKON_INV);
    or TI_OR_GVC_D_D (NOT_TCHKON_OR_GVC_D_D, GVC_D_D, TCHKON_INV);

`endif


specify

      ( CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      ( CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      ( PREZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      ( PREZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_PREZ_PREZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_PREZ_PREZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_D_D != 1 , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge PREZ &&& NOT_TCHKON_OR_Q != 1  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.3 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module DTP23 (CLK , D, PREZ, Q ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input PREZ;
   output Q;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_PREZ_PREZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_pudp   TI_LACTHP_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVC_PREZ_PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_PREZ_PREZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_pudp   TI_LACTHP_UDP2 ( FNET2, D, IINVnet1, PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP3 ( BFONET1, FNET2, CLK, PREZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;



`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_Q_NOTEQ_D_PREZ_NOT0_ , Q , GVC_D_D , 1'bx , 1'b1 , 1'b1 , GVC_PREZ_PREZ ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_PREZ;
    wire TCHKON_AND_GVC_PREZ_PREZ;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_;

    and TI_AND_PREZ (TCHKON_AND_PREZ, PREZ, TCHKON_NET);
    and TI_AND_GVC_PREZ_PREZ (TCHKON_AND_GVC_PREZ_PREZ, GVC_PREZ_PREZ, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_, GVC_Q_NOTEQ_D_PREZ_NOT0_, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_Q;
    wire NOT_TCHKON_OR_D;
    wire NOT_TCHKON_OR_GVC_D_D;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_Q (NOT_TCHKON_OR_Q, Q, TCHKON_INV);
    or TI_OR_D (NOT_TCHKON_OR_D, D, TCHKON_INV);
    or TI_OR_GVC_D_D (NOT_TCHKON_OR_GVC_D_D, GVC_D_D, TCHKON_INV);

`endif


specify

      (CLK  *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_PREZ_PREZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_PREZ_PREZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_D_D != 1 , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge PREZ &&& NOT_TCHKON_OR_Q != 1  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  24-Apr-2000 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module DTP24 (CLK , D, PREZ,  QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input PREZ;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_PREZ_PREZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_pudp   TI_LACTHP_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVC_PREZ_PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_PREZ_PREZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_pudp   TI_LACTHP_UDP2 ( FNET2, D, IINVnet1, PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP3 ( BFONET1, FNET2, CLK, PREZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly


          not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

          not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    not     TI_NOT_PRIM10 (Q, QZ);
    cons_udp TI_COND0 ( GVC_Q_NOTEQ_D_PREZ_NOT0_ , Q , GVC_D_D , 1'bx , 1'b1 , 1'b1 , GVC_PREZ_PREZ ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_PREZ;
    wire TCHKON_AND_GVC_PREZ_PREZ;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_;

    and TI_AND_PREZ (TCHKON_AND_PREZ, PREZ, TCHKON_NET);
    and TI_AND_GVC_PREZ_PREZ (TCHKON_AND_GVC_PREZ_PREZ, GVC_PREZ_PREZ, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_, GVC_Q_NOTEQ_D_PREZ_NOT0_, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_Q;
    wire NOT_TCHKON_OR_D;
    wire NOT_TCHKON_OR_GVC_D_D;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_Q (NOT_TCHKON_OR_Q, Q, TCHKON_INV);
    or TI_OR_D (NOT_TCHKON_OR_D, D, TCHKON_INV);
    or TI_OR_GVC_D_D (NOT_TCHKON_OR_GVC_D_D, GVC_D_D, TCHKON_INV);

`endif


specify

      (CLK  *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_PREZ_PREZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_PREZ_PREZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_D_D != 1 , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge PREZ &&& NOT_TCHKON_OR_Q != 1  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  24-Apr-2000 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module DTP40 (CLK , D, PREZ, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input PREZ;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_PREZ_PREZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_pudp   TI_LACTHP_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVC_PREZ_PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_PREZ_PREZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_pudp   TI_LACTHP_UDP2 ( FNET2, D, IINVnet1, PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP3 ( BFONET1, FNET2, CLK, PREZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_Q_NOTEQ_D_PREZ_NOT0_ , Q , GVC_D_D , 1'bx , 1'b1 , 1'b1 , GVC_PREZ_PREZ ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_PREZ;
    wire TCHKON_AND_GVC_PREZ_PREZ;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_;

    and TI_AND_PREZ (TCHKON_AND_PREZ, PREZ, TCHKON_NET);
    and TI_AND_GVC_PREZ_PREZ (TCHKON_AND_GVC_PREZ_PREZ, GVC_PREZ_PREZ, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_, GVC_Q_NOTEQ_D_PREZ_NOT0_, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_Q;
    wire NOT_TCHKON_OR_D;
    wire NOT_TCHKON_OR_GVC_D_D;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_Q (NOT_TCHKON_OR_Q, Q, TCHKON_INV);
    or TI_OR_D (NOT_TCHKON_OR_D, D, TCHKON_INV);
    or TI_OR_GVC_D_D (NOT_TCHKON_OR_GVC_D_D, GVC_D_D, TCHKON_INV);

`endif


specify

      ( CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      ( CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      ( PREZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      ( PREZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_PREZ_PREZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_PREZ_PREZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_D_D != 1 , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge PREZ &&& NOT_TCHKON_OR_Q != 1  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.3 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module DTP43 (CLK , D, PREZ, Q ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input PREZ;
   output Q;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_PREZ_PREZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_pudp   TI_LACTHP_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVC_PREZ_PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_PREZ_PREZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_pudp   TI_LACTHP_UDP2 ( FNET2, D, IINVnet1, PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP3 ( BFONET1, FNET2, CLK, PREZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;



`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_Q_NOTEQ_D_PREZ_NOT0_ , Q , GVC_D_D , 1'bx , 1'b1 , 1'b1 , GVC_PREZ_PREZ ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_PREZ;
    wire TCHKON_AND_GVC_PREZ_PREZ;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_;

    and TI_AND_PREZ (TCHKON_AND_PREZ, PREZ, TCHKON_NET);
    and TI_AND_GVC_PREZ_PREZ (TCHKON_AND_GVC_PREZ_PREZ, GVC_PREZ_PREZ, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_, GVC_Q_NOTEQ_D_PREZ_NOT0_, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_Q;
    wire NOT_TCHKON_OR_D;
    wire NOT_TCHKON_OR_GVC_D_D;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_Q (NOT_TCHKON_OR_Q, Q, TCHKON_INV);
    or TI_OR_D (NOT_TCHKON_OR_D, D, TCHKON_INV);
    or TI_OR_GVC_D_D (NOT_TCHKON_OR_GVC_D_D, GVC_D_D, TCHKON_INV);

`endif


specify

      (CLK  *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_PREZ_PREZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_PREZ_PREZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_D_D != 1 , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge PREZ &&& NOT_TCHKON_OR_Q != 1  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  24-Apr-2000 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module DTP44 (CLK , D, PREZ,  QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input PREZ;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_PREZ_PREZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_pudp   TI_LACTHP_UDP0 ( FNET2, GVC_D_D, IINVnet1, GVC_PREZ_PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_PREZ_PREZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_pudp   TI_LACTHP_UDP2 ( FNET2, D, IINVnet1, PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP3 ( BFONET1, FNET2, CLK, PREZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly


          not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

          not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    not     TI_NOT_PRIM10 (Q, QZ);
    cons_udp TI_COND0 ( GVC_Q_NOTEQ_D_PREZ_NOT0_ , Q , GVC_D_D , 1'bx , 1'b1 , 1'b1 , GVC_PREZ_PREZ ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_PREZ;
    wire TCHKON_AND_GVC_PREZ_PREZ;
    wire TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_;

    and TI_AND_PREZ (TCHKON_AND_PREZ, PREZ, TCHKON_NET);
    and TI_AND_GVC_PREZ_PREZ (TCHKON_AND_GVC_PREZ_PREZ, GVC_PREZ_PREZ, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_, GVC_Q_NOTEQ_D_PREZ_NOT0_, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_Q;
    wire NOT_TCHKON_OR_D;
    wire NOT_TCHKON_OR_GVC_D_D;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_Q (NOT_TCHKON_OR_Q, Q, TCHKON_INV);
    or TI_OR_D (NOT_TCHKON_OR_D, D, TCHKON_INV);
    or TI_OR_GVC_D_D (NOT_TCHKON_OR_GVC_D_D, GVC_D_D, TCHKON_INV);

`endif


specify

      (CLK  *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_PREZ_PREZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_PREZ_PREZ != 0 , GVC_CLK_CLK, GVC_D_D ); 
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_D_D != 1 , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge PREZ &&& NOT_TCHKON_OR_Q != 1  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  24-Apr-2000 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module EN210 ( A, B, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input A ;
        input B ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           xnor #0 TI_XNOR_PRIM0 ( Y, A, B ) ;

      `ifdef TI_functiononly
`else
      specify
             if (!B)
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if (B)
                ( A => Y ) = ( 0.0100, 0.0100 ) ;

             if (!A)
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if (A)
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify



`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module EN220 ( A, B, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input A ;
        input B ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           xnor #0 TI_XNOR_PRIM0 ( Y, A, B ) ;

      `ifdef TI_functiononly
`else
      specify
             if (!B)
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if (B)
                ( A => Y ) = ( 0.0100, 0.0100 ) ;

             if (!A)
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if (A)
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify



`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module EN240 ( A, B, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input A ;
        input B ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           xnor #0 TI_XNOR_PRIM0 ( Y, A, B ) ;

      `ifdef TI_functiononly
`else
      specify
             if (!B)
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if (B)
                ( A => Y ) = ( 0.0100, 0.0100 ) ;

             if (!A)
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if (A)
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify



`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module EN310 ( A, B, C, Y ) ;

 // Verilog Port Declaration section
       output Y ;
        input A ;
        input B ;
        input C ;

    `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           xnor #0 TI_XNOR_PRIM0 ( Y, A, B, C ) ;

     `ifdef TI_functiononly
`else
       specify
             if(!B && !C)
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if(!B && C)
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if(B && !C)
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if(B && C)
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             
             if(!A && !C)
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if(!A && C)
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if(A && !C)
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if(A && C)
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             
             if(!A && !B)
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if(!A && B)
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if(A && !B)
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if(A && B)
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module EN320 ( A, B, C, Y ) ;

 // Verilog Port Declaration section
       output Y ;
        input A ;
        input B ;
        input C ;

    `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           xnor #0 TI_XNOR_PRIM0 ( Y, A, B, C ) ;

     `ifdef TI_functiononly
`else
       specify
             if(!B && !C)
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if(!B && C)
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if(B && !C)
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if(B && C)
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             
             if(!A && !C)
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if(!A && C)
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if(A && !C)
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if(A && C)
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             
             if(!A && !B)
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if(!A && B)
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if(A && !B)
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if(A && B)
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module EN340 ( A, B, C, Y ) ;

 // Verilog Port Declaration section
       output Y ;
        input A ;
        input B ;
        input C ;

    `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           xnor #0 TI_XNOR_PRIM0 ( Y, A, B, C ) ;

     `ifdef TI_functiononly
`else
       specify
             if(!B && !C)
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if(!B && C)
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if(B && !C)
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if(B && C)
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             
             if(!A && !C)
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if(!A && C)
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if(A && !C)
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if(A && C)
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             
             if(!A && !B)
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if(!A && B)
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if(A && !B)
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if(A && B)
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module EX210 ( A, B, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input A ;
        input B ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

           xor #0 TI_XOR_PRIM0 ( Y, A, B ) ;
    `ifdef TI_functiononly
`else

        specify
             if (!B)
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if (B)
                ( A => Y ) = ( 0.0100, 0.0100 ) ;

             if (!A)
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if (A)
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module EX220 ( A, B, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input A ;
        input B ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

           xor #0 TI_XOR_PRIM0 ( Y, A, B ) ;
    `ifdef TI_functiononly
`else

        specify
             if (!B)
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if (B)
                ( A => Y ) = ( 0.0100, 0.0100 ) ;

             if (!A)
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if (A)
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module EX240 ( A, B, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input A ;
        input B ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

           xor #0 TI_XOR_PRIM0 ( Y, A, B ) ;
    `ifdef TI_functiononly
`else

        specify
             if (!B)
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if (B)
                ( A => Y ) = ( 0.0100, 0.0100 ) ;

             if (!A)
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if (A)
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module EX310 ( A, B, C, Y ) ;

   // Verilog Port Declaration section
        output Y ;
        input A ;
        input B ;
        input C ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           xor #0 TI_XOR_PRIM0 ( Y, A, B, C ) ;

     `ifdef TI_functiononly
`else
       specify
             if (!B && !C )
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if (!B && C )
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if (B && !C )
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if (B && C )
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;

             if (!A && !C )
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if (A && C )
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if (A && !C )
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if (!A && C )
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;

             if (!A && !B )
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if (A && !B )
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if (A && B )
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if (!A && B )
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module EX320 ( A, B, C, Y ) ;

   // Verilog Port Declaration section
        output Y ;
        input A ;
        input B ;
        input C ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           xor #0 TI_XOR_PRIM0 ( Y, A, B, C ) ;

     `ifdef TI_functiononly
`else
       specify
             if (!B && !C )
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if (!B && C )
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if (B && !C )
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if (B && C )
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;

             if (!A && !C )
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if (A && C )
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if (A && !C )
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if (!A && C )
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;

             if (!A && !B )
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if (A && !B )
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if (A && B )
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if (!A && B )
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module EX340 ( A, B, C, Y ) ;

   // Verilog Port Declaration section
        output Y ;
        input A ;
        input B ;
        input C ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           xor #0 TI_XOR_PRIM0 ( Y, A, B, C ) ;

     `ifdef TI_functiononly
`else
       specify
             if (!B && !C )
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if (!B && C )
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if (B && !C )
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;
             if (B && C )
                  ( A => Y ) = ( 0.0100, 0.0100 ) ;

             if (!A && !C )
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if (A && C )
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if (A && !C )
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;
             if (!A && C )
                  ( B => Y ) = ( 0.0100, 0.0100 ) ;

             if (!A && !B )
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if (A && !B )
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if (A && B )
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
             if (!A && B )
                  ( C => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module FA320P ( A, B, CI, CO, S ) ;

// Verilog Port Declaration section
        output CO ;
        output S ;
        input A ;
        input B ;
        input CI ;
        
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
        and TI_AND_PRIM0 ( NODE1, A, B ) ;
        and TI_AND_PRIM1 ( NODE2, B, CI ) ;
        and TI_AND_PRIM2 ( NODE3, CI, A ) ;
        or #0 TI_OR_PRIM0 ( CO, NODE1, NODE2, NODE3 ) ;
        xor #0 TI_XOR_PRIM0 ( S, A, B, CI ) ;

    `ifdef TI_functiononly
`else
        specify
             if (B && !CI )
                  ( A => CO ) = ( 0.0100, 0.0100 ) ;
             if (!B && CI )
                  ( A => CO ) = ( 0.0100, 0.0100 ) ;

             if (A && !CI )
                  ( B => CO ) = ( 0.0100, 0.0100 ) ;
             if (!A && CI )
                  ( B => CO ) = ( 0.0100, 0.0100 ) ;

             if (A && !B )
                  ( CI => CO ) = ( 0.0100, 0.0100 ) ;
             if (!A && B )
                  ( CI => CO ) = ( 0.0100, 0.0100 ) ;

             if (!B && !CI )
                  ( A => S ) = ( 0.0100, 0.0100 ) ;
             if (!B && CI )
                  ( A => S ) = ( 0.0100, 0.0100 ) ;
             if (B && !CI )
                  ( A => S ) = ( 0.0100, 0.0100 ) ;
             if (B && CI )
                  ( A => S ) = ( 0.0100, 0.0100 ) ;

             if (!A && !CI )
                  ( B => S ) = ( 0.0100, 0.0100 ) ;
             if (A && CI )
                  ( B => S ) = ( 0.0100, 0.0100 ) ;
             if (A && !CI )
                  ( B => S ) = ( 0.0100, 0.0100 ) ;
             if (!A && CI )
                  ( B => S ) = ( 0.0100, 0.0100 ) ;

             if (!A && !B )
                  ( CI => S ) = ( 0.0100, 0.0100 ) ;
             if (A && !B )
                  ( CI => S ) = ( 0.0100, 0.0100 ) ;
             if (A && B )
                  ( CI => S ) = ( 0.0100, 0.0100 ) ;
             if (!A && B )
                  ( CI => S ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module FA320 ( A, B, CI, CO, S ) ;

// Verilog Port Declaration section
        output CO ;
        output S ;
        input A ;
        input B ;
        input CI ;
        
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
        and TI_AND_PRIM0 ( NODE1, A, B ) ;
        and TI_AND_PRIM1 ( NODE2, B, CI ) ;
        and TI_AND_PRIM2 ( NODE3, CI, A ) ;
        or #0 TI_OR_PRIM0 ( CO, NODE1, NODE2, NODE3 ) ;
        xor #0 TI_XOR_PRIM0 ( S, A, B, CI ) ;

    `ifdef TI_functiononly
`else
        specify
             if (B && !CI )
                  ( A => CO ) = ( 0.0100, 0.0100 ) ;
             if (!B && CI )
                  ( A => CO ) = ( 0.0100, 0.0100 ) ;

             if (A && !CI )
                  ( B => CO ) = ( 0.0100, 0.0100 ) ;
             if (!A && CI )
                  ( B => CO ) = ( 0.0100, 0.0100 ) ;

             if (A && !B )
                  ( CI => CO ) = ( 0.0100, 0.0100 ) ;
             if (!A && B )
                  ( CI => CO ) = ( 0.0100, 0.0100 ) ;

             if (!B && !CI )
                  ( A => S ) = ( 0.0100, 0.0100 ) ;
             if (!B && CI )
                  ( A => S ) = ( 0.0100, 0.0100 ) ;
             if (B && !CI )
                  ( A => S ) = ( 0.0100, 0.0100 ) ;
             if (B && CI )
                  ( A => S ) = ( 0.0100, 0.0100 ) ;

             if (!A && !CI )
                  ( B => S ) = ( 0.0100, 0.0100 ) ;
             if (A && CI )
                  ( B => S ) = ( 0.0100, 0.0100 ) ;
             if (A && !CI )
                  ( B => S ) = ( 0.0100, 0.0100 ) ;
             if (!A && CI )
                  ( B => S ) = ( 0.0100, 0.0100 ) ;

             if (!A && !B )
                  ( CI => S ) = ( 0.0100, 0.0100 ) ;
             if (A && !B )
                  ( CI => S ) = ( 0.0100, 0.0100 ) ;
             if (A && B )
                  ( CI => S ) = ( 0.0100, 0.0100 ) ;
             if (!A && B )
                  ( CI => S ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module FA340P ( A, B, CI, CO, S ) ;

// Verilog Port Declaration section
        output CO ;
        output S ;
        input A ;
        input B ;
        input CI ;
        
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
        and TI_AND_PRIM0 ( NODE1, A, B ) ;
        and TI_AND_PRIM1 ( NODE2, B, CI ) ;
        and TI_AND_PRIM2 ( NODE3, CI, A ) ;
        or #0 TI_OR_PRIM0 ( CO, NODE1, NODE2, NODE3 ) ;
        xor #0 TI_XOR_PRIM0 ( S, A, B, CI ) ;

    `ifdef TI_functiononly
`else
        specify
             if (B && !CI )
                  ( A => CO ) = ( 0.0100, 0.0100 ) ;
             if (!B && CI )
                  ( A => CO ) = ( 0.0100, 0.0100 ) ;

             if (A && !CI )
                  ( B => CO ) = ( 0.0100, 0.0100 ) ;
             if (!A && CI )
                  ( B => CO ) = ( 0.0100, 0.0100 ) ;

             if (A && !B )
                  ( CI => CO ) = ( 0.0100, 0.0100 ) ;
             if (!A && B )
                  ( CI => CO ) = ( 0.0100, 0.0100 ) ;

             if (!B && !CI )
                  ( A => S ) = ( 0.0100, 0.0100 ) ;
             if (!B && CI )
                  ( A => S ) = ( 0.0100, 0.0100 ) ;
             if (B && !CI )
                  ( A => S ) = ( 0.0100, 0.0100 ) ;
             if (B && CI )
                  ( A => S ) = ( 0.0100, 0.0100 ) ;

             if (!A && !CI )
                  ( B => S ) = ( 0.0100, 0.0100 ) ;
             if (A && CI )
                  ( B => S ) = ( 0.0100, 0.0100 ) ;
             if (A && !CI )
                  ( B => S ) = ( 0.0100, 0.0100 ) ;
             if (!A && CI )
                  ( B => S ) = ( 0.0100, 0.0100 ) ;

             if (!A && !B )
                  ( CI => S ) = ( 0.0100, 0.0100 ) ;
             if (A && !B )
                  ( CI => S ) = ( 0.0100, 0.0100 ) ;
             if (A && B )
                  ( CI => S ) = ( 0.0100, 0.0100 ) ;
             if (!A && B )
                  ( CI => S ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module FA340 ( A, B, CI, CO, S ) ;

// Verilog Port Declaration section
        output CO ;
        output S ;
        input A ;
        input B ;
        input CI ;
        
 `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
        and TI_AND_PRIM0 ( NODE1, A, B ) ;
        and TI_AND_PRIM1 ( NODE2, B, CI ) ;
        and TI_AND_PRIM2 ( NODE3, CI, A ) ;
        or #0 TI_OR_PRIM0 ( CO, NODE1, NODE2, NODE3 ) ;
        xor #0 TI_XOR_PRIM0 ( S, A, B, CI ) ;

    `ifdef TI_functiononly
`else
        specify
             if (B && !CI )
                  ( A => CO ) = ( 0.0100, 0.0100 ) ;
             if (!B && CI )
                  ( A => CO ) = ( 0.0100, 0.0100 ) ;

             if (A && !CI )
                  ( B => CO ) = ( 0.0100, 0.0100 ) ;
             if (!A && CI )
                  ( B => CO ) = ( 0.0100, 0.0100 ) ;

             if (A && !B )
                  ( CI => CO ) = ( 0.0100, 0.0100 ) ;
             if (!A && B )
                  ( CI => CO ) = ( 0.0100, 0.0100 ) ;

             if (!B && !CI )
                  ( A => S ) = ( 0.0100, 0.0100 ) ;
             if (!B && CI )
                  ( A => S ) = ( 0.0100, 0.0100 ) ;
             if (B && !CI )
                  ( A => S ) = ( 0.0100, 0.0100 ) ;
             if (B && CI )
                  ( A => S ) = ( 0.0100, 0.0100 ) ;

             if (!A && !CI )
                  ( B => S ) = ( 0.0100, 0.0100 ) ;
             if (A && CI )
                  ( B => S ) = ( 0.0100, 0.0100 ) ;
             if (A && !CI )
                  ( B => S ) = ( 0.0100, 0.0100 ) ;
             if (!A && CI )
                  ( B => S ) = ( 0.0100, 0.0100 ) ;

             if (!A && !B )
                  ( CI => S ) = ( 0.0100, 0.0100 ) ;
             if (A && !B )
                  ( CI => S ) = ( 0.0100, 0.0100 ) ;
             if (A && B )
                  ( CI => S ) = ( 0.0100, 0.0100 ) ;
             if (!A && B )
                  ( CI => S ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module HA220 ( A, B, CO, S ) ;

// Verilog Port Declaration section
        output CO ;
        output S ;
        input A ;
        input B ;
        
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           and #0 TI_AND_PRIM0 ( CO, A, B ) ;
           xor #0 TI_XOR_PRIM0 ( S, A, B ) ;
        
    `ifdef TI_functiononly
`else
    specify
                ( A *> CO ) = ( 0.0100, 0.0100 ) ;
                ( B *> CO ) = ( 0.0100, 0.0100 ) ;

             if (!B )
                  ( A *> S ) = ( 0.0100, 0.0100 ) ;
             if (B )
                  ( A *> S ) = ( 0.0100, 0.0100 ) ;

             if (!A )
                  ( B *> S ) = ( 0.0100, 0.0100 ) ;
             if (A )
                  ( B *> S ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module HA221 ( A, B, CO, S ) ;

   // Verilog Port Declaration section
        output CO ;
        output S ;
        input A ;
        input B ;
   `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

     
           or #0 TI_OR_PRIM0 ( CO, A, B ) ;
           xnor #0 TI_XNOR_PRIM0 ( S, A, B ) ;
        
`ifdef TI_functiononly
`else

        specify
                ( A *> CO ) = ( 0.0100, 0.0100 ) ;
                ( B *> CO ) = ( 0.0100, 0.0100 ) ;

             if (!B )
                  ( A *> S ) = ( 0.0100, 0.0100 ) ;
             if (B )
                  ( A *> S ) = ( 0.0100, 0.0100 ) ;

             if (!A )
                  ( B *> S ) = ( 0.0100, 0.0100 ) ;
             if (A )
                  ( B *> S ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module IV110 ( A, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           not #0 TI_NOT_PRIM0 ( Y, A ) ;
`ifdef TI_functiononly
`else


        specify
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module IV120 ( A, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           not #0 TI_NOT_PRIM0 ( Y, A ) ;
`ifdef TI_functiononly
`else


        specify
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module IV130 ( A, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           not #0 TI_NOT_PRIM0 ( Y, A ) ;
`ifdef TI_functiononly
`else


        specify
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module IV140 ( A, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           not #0 TI_NOT_PRIM0 ( Y, A ) ;
`ifdef TI_functiononly
`else


        specify
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module IV180 ( A, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           not #0 TI_NOT_PRIM0 ( Y, A ) ;
`ifdef TI_functiononly
`else


        specify
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module IV190 ( A, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           not #0 TI_NOT_PRIM0 ( Y, A ) ;
`ifdef TI_functiononly
`else


        specify
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module IV1G0 ( A, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           not #0 TI_NOT_PRIM0 ( Y, A ) ;
`ifdef TI_functiononly
`else


        specify
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module IV1W0 ( A, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
           not #0 TI_NOT_PRIM0 ( Y, A ) ;
`ifdef TI_functiononly
`else


        specify
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module IV240 ( A, G, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A ;
        input G ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        notif1 #0 TI_NOTIF1_PRIM0( Y, A, G) ;

`ifdef TI_functiononly
`else
        specify
                ( G => Y ) = ( 0.0100, 0.0100, 0.0100, 0.0100, 0.0100, 0.0100 ) ;
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module IV280 ( A, G, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A ;
        input G ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        notif1 #0 TI_NOTIF1_PRIM0( Y, A, G) ;

`ifdef TI_functiononly
`else
        specify
                ( G => Y ) = ( 0.0100, 0.0100, 0.0100, 0.0100, 0.0100, 0.0100 ) ;
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module IV2G0 ( A, G, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A ;
        input G ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        notif1 #0 TI_NOTIF1_PRIM0( Y, A, G) ;

`ifdef TI_functiononly
`else
        specify
                ( G => Y ) = ( 0.0100, 0.0100, 0.0100, 0.0100, 0.0100, 0.0100 ) ;
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module IV2P0 ( A, G, Y ) ;
// Verilog Port Declaration section

        output Y ;
        input A ;
        input G ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        notif1 #0 TI_NOTIF1_PRIM0( Y, A, G) ;

`ifdef TI_functiononly
`else
        specify
                ( G => Y ) = ( 0.0100, 0.0100, 0.0100, 0.0100, 0.0100, 0.0100 ) ;
                ( A => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly    
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module LAB20 (CLRZ, D, ENZ, PREZ, Q, QZ ) ;

// Verilog Port Declaration section

   input CLRZ;
   input D;
   input ENZ;
   input PREZ;
   output Q;
   output QZ;

`ifdef TI_verilog    
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
    parameter Xon = 1;
    wire GVCnotifier1;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;

// Xon controlability

   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_ENZ_ENZ ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ,  GVC_PREZ_PREZ  ; 

           not      ( NOT_GVC_ENZ_ENZ, GVC_ENZ_ENZ ) ;
         laudp_msl   TI_LATCH_UDP0 ( BFONET1, GVC_D_D, NOT_GVC_ENZ_ENZ, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier1 ) ;
       laqzudp_msl   TI_LAQZ_UDP0 ( BFONET2, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, BFONET1 ) ;


`else
 
           not      ( NOT_ENZ, ENZ ) ;
         laudp_msl   TI_LATCH_UDP1 ( BFONET1, D, NOT_ENZ, CLRZ, PREZ, GVCnotifier1 ) ;
       laqzudp_msl   TI_LAQZ_UDP1 ( BFONET2, CLRZ, PREZ, BFONET1 ) ;


`endif

`ifdef TI_functiononly
 
          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          buf #1 TI_BUF_PRIM1 ( QZ, BFONET2 ) ;


`else

          buf  TI_BUF_PRIM2 ( Q, BFONET1 ) ;
          buf  TI_BUF_PRIM3 ( QZ, BFONET2 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_CLRZ_NOT0_PREZ_NOT0_ , 1'b0 , 1'b1 , 1'bx , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOT0_PREZ_NOT0_ , GVC_D_D , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_D_NOT1_CLRZ_NOT0_ , GVC_D_D , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_D_NOTEQ_Q_CLRZ_NOT0_PREZ_NOT0 , GVC_D_D , Q , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND4 ( GVC_Q_NOT0_PREZ_NOT0_ , Q , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND5 ( GVC_Q_NOT1_CLRZ_NOT0_ , Q , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly


specify
    $recovery(posedge PREZ ,posedge CLRZ &&& ( ENZ != 0 ) ,1,GVCnotifier1_zd );
endspecify

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0_PREZ_NOT0;
    wire TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_;

    and TI_AND_GVC_D_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_, GVC_D_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_, GVC_Q_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_, GVC_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0_PREZ_NOT0 (TCHKON_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0_PREZ_NOT0, GVC_D_NOTEQ_Q_CLRZ_NOT0_PREZ_NOT0, TCHKON_NET);
    and TI_AND_GVC_D_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_, GVC_D_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_, GVC_Q_NOT1_CLRZ_NOT0_, TCHKON_NET);

    wire TCHKON_AND_GVC_ENZ_ENZ;
    wire TCHKON_AND_ENZ;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    and TI_AND_GVC_ENZ_ENZ (TCHKON_AND_GVC_ENZ_ENZ, GVC_ENZ_ENZ, TCHKON_NET);
    and TI_AND_ENZ (TCHKON_AND_ENZ, ENZ, TCHKON_NET);

`endif


specify
      (ENZ    *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (ENZ    *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ   *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ   *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (D      *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (D      *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ   *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ   *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge ENZ,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ != 0 ) , GVC_ENZ_ENZ, GVC_D_D ); 
   $setuphold(posedge ENZ,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_CLRZ_NOT0_PREZ_NOT0_ != 0 ) , GVC_ENZ_ENZ, GVC_D_D ); 
   $recrem(posedge CLRZ,  posedge ENZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_D_NOT0_PREZ_NOT0_ != 0 ) , GVC_CLRZ_CLRZ , GVC_ENZ_ENZ);
   $recrem(posedge PREZ,  posedge ENZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_D_NOT1_CLRZ_NOT0_ != 0 ) , GVC_PREZ_PREZ , GVC_ENZ_ENZ);
   $setuphold(posedge PREZ, posedge CLRZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_ENZ_ENZ != 0 ), GVC_PREZ_PREZ, GVC_CLRZ_CLRZ ); 
   $setuphold(posedge CLRZ, posedge PREZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_ENZ_ENZ != 0 ), GVC_CLRZ_CLRZ, GVC_PREZ_PREZ ); 
   $width(negedge ENZ  &&& ( TCHKON_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0_PREZ_NOT0 != 0 )  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ  &&& ( TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_ != 0 )  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge PREZ  &&& ( TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_ != 0 )  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

//#------------------------------------------------------------
//# Revision History
//# Last Modified on:  Wed Aug 17 2005
//# Modifications: 
//# a) Verilog Port Declaration section:
//#    Change in the Port order, in sync with module defination
//#------------------------------------------------------------

// Revision history:
// ----------------

//v1.1 09-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module LAC20 (CLRZ , ENZ, D, Q, QZ ) ;

// Verilog Port Declaration section

   input CLRZ;
   input ENZ;
   input D;
   output Q;
   output QZ;

`ifdef TETRAMAX

  _DLAT L1 ( 1'b0,!CLRZ,!ENZ,D,QINT);
  _AND  A1 ( CLRZ, QINT, Q);
  _INV  I1 ( QINT, QZINT);
  _OR   A2 ( QZINT, !CLRZ, QZ);

`else

`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_ENZ_ENZ ,  GVC_D_D  ,  GVC_CLRZ_CLRZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_ENZ_ENZ ) ;
       la_cudp   TI_LACTHC_UDP0 ( BFONET1, GVC_D_D, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, ENZ ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, D, IINVnet1, CLRZ, GVCnotifier1 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM2 ( QZ, BFONET1 );


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM3 ( QZ, BFONET1 );

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_D_NOTEQ_Q_CLRZ_NOT0 , GVC_D_D , Q , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_CLRZ_CLRZ;
    wire TCHKON_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0;
    wire TCHKON_AND_Q;
    wire TCHKON_AND_D;
    wire TCHKON_AND_GVC_D_D;
    wire TCHKON_AND_CLRZ;

    and TI_AND_GVC_CLRZ_CLRZ (TCHKON_AND_GVC_CLRZ_CLRZ, GVC_CLRZ_CLRZ, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0 (TCHKON_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0, GVC_D_NOTEQ_Q_CLRZ_NOT0, TCHKON_NET);
    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_D (TCHKON_AND_D, D, TCHKON_NET);
    and TI_AND_GVC_D_D (TCHKON_AND_GVC_D_D, GVC_D_D, TCHKON_NET);
    and TI_AND_CLRZ (TCHKON_AND_CLRZ, CLRZ, TCHKON_NET);

`endif


specify

      (D    *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (ENZ   *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (D    *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (ENZ   *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge ENZ,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_ENZ_ENZ, GVC_D_D ); 
   $setuphold(posedge ENZ,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_CLRZ_CLRZ != 0 , GVC_ENZ_ENZ, GVC_D_D ); 
   $recrem(posedge CLRZ,  posedge ENZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_D != 0 , GVC_CLRZ_CLRZ , GVC_ENZ_ENZ);
   $width(negedge CLRZ &&& TCHKON_AND_Q != 0  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge ENZ  &&& TCHKON_AND_GVC_D_NOTEQ_Q_CLRZ_NOT0 != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

`endif // ifdef TETRAMAX
endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.5 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.

// v1.4  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.3  05-Sep-2001 Removed the Copyright block
// v1.2  11-Apr-2000 Updated for Tetramax support
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2002 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

`resetall

`ifdef TI_functiononly
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif
primitive la_cudp(q, d, c, clr, nt);

input d, c, clr, nt;
output q;
reg q;

table
//	d	c  clr  nt  :q:  q;

	?	?  (?0)	?   :?:	 0;
	*	?   0	?   :?:	 0;
	?	*   0	?   :?:	 0;

        (?0)    ?   ?	?   :0:  0;
    	0  	*   ?   ?   :0:	 0;
    	0       ?   *   ?   :0:	 0;

	?      (?0) 1	?   :?:	 -;
	?	0 (?1)  ?   :?:	 -;
	*	0   1   ?   :?:	 -;

//reduction of pessimism
  	(?0)	1  ?    ?   :?:	 0;
	0 (?1)  ?	?   :?:	 0;
	0	1  *    ?   :?:	 0;

  	(?1)  1	1	?   :?:  1;
	1 (?1)  1	?   :?:	 1;
	1	1 (?1)  ?   :?:	 1;

   	(?1) ?   1	?   :1:  1;
    	1   ? (?1)	?   :1:	 1;
    	1   *   1	?   :1:	 1;

	? (?0)	x	?   :0:  0;
	?	0 (?x)  ?   :0:	 0;
	*	0   x   ?   :0:	 0;

	?	?	?   *   :?:  x;

endtable
endprimitive 

// Revision history:
// ----------------
// v1.2  08-Jun-1999  Changing 10ps to 1ps
// v1.1  17-Mar-1999 24 date and time created 99/03/17 17
// v1.2  08-Jun-1999  Changing 10ps to 1ps
// v1.1  17-Mar-1999 24 date and time created 99/03/17 17
// 19 Dec 2006 : Sharavathi : changed the timescale for functiononly option to 
//                            1ns/1ps
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module LAN20 (D, ENZ , Q, QZ ) ;

// Verilog Port Declaration section
   input D;
   input ENZ;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_ENZ_ENZ ,  GVC_D_D  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_ENZ_ENZ ) ;
       la_nudp   TI_LACTHN_UDP0 ( BFONET1, GVC_D_D, IINVnet1, GVCnotifier1 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, ENZ ) ;
       la_nudp   TI_LACTHN_UDP1 ( BFONET1, D, IINVnet1, GVCnotifier1 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_D_NOTEQ_Q , GVC_D_D , Q , 1'b0 , 1'b1 , 1'b1 , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_D_NOTEQ_Q;

    and TI_AND_GVC_D_NOTEQ_Q (TCHKON_AND_GVC_D_NOTEQ_Q, GVC_D_NOTEQ_Q, TCHKON_NET);

`endif


specify

      (D  *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (D  *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (ENZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (ENZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge ENZ &&& (TCHKON_NET != 0) ,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_ENZ_ENZ, GVC_D_D ); 
   $setuphold(posedge ENZ &&& (TCHKON_NET != 0) ,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,, GVC_ENZ_ENZ, GVC_D_D ); 
   $width(negedge ENZ  &&& TCHKON_AND_GVC_D_NOTEQ_Q != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.5 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.4  17-Aug-2005 Verilog Port Declaration section:Change in the Port order,
//                   in sync with module defination
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2002 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

`resetall

`ifdef TI_functiononly
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif
primitive la_nudp(q, d, c, nt);

input d, c, nt;
output q;
reg q;

table
//	d   c     nt   :q:  q;

	?  (?0)   ?    :?:  -;
	*   0	  ?    :?:  -;

//reduction of pessimism

       (?0) 1	  ?    :?:  0;
	0  (?1)   ?    :?:  0;

       (?1) 1	  ?    :?:  1;
	1  (?1)   ?    :?:  1;

       (?1) ?     ?    :1:  1;
        1   *     ?    :1:  1;

       (?0) ?	  ?    :0:  0;
        0   *     ?    :0:  0;

	?   ?	  *    :?:  x;

// not  pz  cz  c  cih  d  sd  tc : q0 : q TSCZ  MSt   St   MSt    Q   QZ   SQ

//if PREZ = 0 and CLRZ = 1;
//   ?    0   1   1   ?   0  0   1  : ?  : 0 ;

   // when TMC is X
//   ?    0   1   1   ?   0  0   X  0  ?  ?  X  X 0 X;

endtable
endprimitive 
// Revision history:
// ----------------
// v1.2  08-Jun-1999  Changing 10ps to 1ps
// v1.1  17-Mar-1999 24 date and time created 99/03/17 17
// v1.2  08-Jun-1999  Changing 10ps to 1ps
// v1.1  17-Mar-1999 24 date and time created 99/03/17 17
// 19 Dec 2006 : Sharavathi : changed the timescale for functiononly option to 
//                            1ns/1ps
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module LAP20 (D, ENZ, PREZ, Q, QZ  ) ;

// Verilog Port Declaration section
   input D;
   input ENZ;
   input PREZ;
   output Q;
   output QZ;

`ifdef TI_verilog    
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
    parameter Xon = 1;
    wire GVCnotifier1;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;

// Xon controlability

   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_ENZ_ENZ ,  GVC_D_D  ,    GVC_PREZ_PREZ  ; 

           not   TI_NOT_PRIM0 ( IINVnet1, GVC_ENZ_ENZ ) ;
       la_pudp   TI_LACTHC_UDP0 ( BFONET1, GVC_D_D, IINVnet1, GVC_PREZ_PREZ, GVCnotifier1 ) ;


`else

           not   TI_NOT_PRIM1 ( IINVnet1, ENZ ) ;
       la_pudp   TI_LACTHC_UDP1 ( BFONET1, D, IINVnet1, PREZ, GVCnotifier1 ) ;


`endif


`ifdef TI_functiononly
 
          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_BUF_PRIM1 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM2 ( Q, BFONET1 ) ;
          not  TI_BUF_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_D_NOTEQ_Q_PREZ_NOT0_ , GVC_D_D , Q , 1'b0 , 1'b1 , 1'b1 , GVC_PREZ_PREZ ) ;

`endif


`ifdef TI_functiononly


`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_D_NOTEQ_Q_PREZ_NOT0_;
    wire TCHKON_AND_GVC_PREZ_PREZ;
    wire TCHKON_AND_PREZ;

    and TI_AND_GVC_D_NOTEQ_Q_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_Q_PREZ_NOT0_, GVC_D_NOTEQ_Q_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_PREZ_PREZ (TCHKON_AND_GVC_PREZ_PREZ, GVC_PREZ_PREZ, TCHKON_NET);
    and TI_AND_PREZ (TCHKON_AND_PREZ, PREZ, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_Q;
    wire NOT_TCHKON_OR_D;
    wire NOT_TCHKON_OR_GVC_D_D;
    
    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_Q (NOT_TCHKON_OR_Q, Q, TCHKON_INV);
    or TI_OR_D (NOT_TCHKON_OR_D, D, TCHKON_INV);
    or TI_OR_GVC_D_D (NOT_TCHKON_OR_GVC_D_D, GVC_D_D, TCHKON_INV);
    
`endif


specify
      (ENZ    *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (ENZ    *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (D      *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (D      *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ   *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ   *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge ENZ,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_PREZ_PREZ != 0 ), GVC_ENZ_ENZ, GVC_D_D ); 
   $setuphold(posedge ENZ,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_PREZ_PREZ != 0 ), GVC_ENZ_ENZ, GVC_D_D ); 
   $recrem(posedge PREZ,  posedge ENZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( NOT_TCHKON_OR_GVC_D_D != 1 ), GVC_PREZ_PREZ , GVC_ENZ_ENZ);
   $width(negedge PREZ &&& ( NOT_TCHKON_OR_Q != 1 ) ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge ENZ  &&& ( TCHKON_AND_GVC_D_NOTEQ_Q_PREZ_NOT0_ != 0 )  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 


`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

//#------------------------------------------------------------
//# Revision History
//# Last Modified on:  Wed Aug 17 2005
//# v1.5 Verilog Port Declaration section: Change in the Port order,
//#      in sync with module defination
//#------------------------------------------------------------

// Revision history:
// ----------------

//v1.1 09-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2002 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

`resetall

`ifdef TI_functiononly
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif
primitive la_pudp(q, d, c, pre, nt);

input d, c,  pre, nt;
output q;
reg q;

table
//	d	c  pre  nt  :q:  q;

	*	?	0   ?   :?:	 1;//
	?	*	0   ?   :?:  1;//
	?	?  (?0) ?   :?:  1;//

   (?1) ?   ?   ?   :1:	 1;
    1   *   ?   ?   :1:  1;
    1   ?   *   ?   :1:  1;

	? (?0)  1   ?   :?:  -;
	?	0  (?1) ?   :?:  -;
	*	0   1   ?   :?:  -;

//reduction of pessimism
  (?0)	1	1   ?   :?:	 0;
	0 (?1)  1   ?   :?:  0;
	0	1  (?1) ?   :?:  0;

  (?1)  1	?   ?   :?:  1;
	1 (?1)  ?   ?   :?:  1;
	1	1   *   ?   :?:	 1;

  (?0)  ?	1   ?   :0:  0;
    0   ?  (?1) ?   :0:	 0;
    0  	*   1   ?   :0:  0;

	? (?0)	x   ?   :1:  1;
	?	0  (?x) ?   :1:  1;
	*	0   x   ?   :1:  1; 

	?	?	?   *   :?:  x;

endtable
endprimitive

// Revision history:
// ----------------
// v1.2  08-Jun-1999  Changing 10ps to 1ps
// v1.1  17-Mar-1999 24 date and time created 99/03/17 17
// v1.2  08-Jun-1999  Changing 10ps to 1ps
// v1.1  17-Mar-1999 24 date and time created 99/03/17 17
// 19 Dec 2006 : Sharavathi : changed the timescale for functiononly option to 
//                            1ns/1ps 
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
`resetall
`ifdef TI_functiononly
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

primitive laqzudp_msl
`protect
(qz, clrz, prez, q);
input clrz, prez, q;
output qz;
table
// clrz prez q qz
    0    ?   ? :1;
    ?    1   0 :1;
    1    0   ? :0;
    1    ?   1 :0;
endtable
`endprotect
endprimitive 

// 19 Dec 2006 : Sharavathi : changed the timescale for functiononly option to 
//                            1ns/1ps

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed

`resetall

`ifdef TI_functiononly
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

primitive laudp_msl
`protect
(q, d, c, clr, pre, nt);

input d, c, clr, pre, nt;
output q;
reg q;

table
//  d   c  clr pre nt  :q:  q;

    ?   ?  (?0) ?  ?   :?:  0;
    *   ?   0   ?  ?   :?:  0;
    ?   *   0   ?  ?   :?:  0;
    ?   ?   0   *  ?   :?:  0;

    ?   ?   1 (?0) ?   :?:  1;
    *   ?   1   0  ?   :?:  1;
    ?   *   1   0  ?   :?:  1;
    ?   ?  (?1) 0  ?   :?:  1;

   (?1) ?   1   ?  ?   :1:  1;
    1   *   1   ?  ?   :1:  1;
    1   ? (?1)  ?  ?   :1:  1;
    1   ?   1   *  ?   :1:  1;

  (?0)  ?   ?   1  ?   :0:  0;
    0   *   ?   1  ?   :0:  0;
    0   ?   *   1  ?   :0:  0;
    0   ?   ? (?1) ?   :0:  0;

    ? (?0)  1   1  ?   :?:  -;
    ?   0 (?1)  1  ?   :?:  -;
    ?   0   1 (?1) ?   :?:  -;
    *   0   1   1  ?   :?:  -;
//reduction of pessimism
  (?0)  1   ?   1  ?   :?:  0;
    0 (?1)  ?   1  ?   :?:  0;
    0   1   ? (?1) ?   :?:  0;
    0   1   *   1  ?   :?:  0;

  (?1)  1   1   ?  ?   :?:  1;
    1 (?1)  1   ?  ?   :?:  1;
    1   1 (?1)  ?  ?   :?:  1;
    1   1   1   *  ?   :?:  1;

    ? (?0)  x   1  ?   :0:  0;
    ?   0 (?x)  1  ?   :0:  0;
    ?   0   x (?1) ?   :0:  0;
    *   0   x   1  ?   :0:  0;

    ? (?0)  1   x  ?   :1:  1;
    ?   0  (?1) x  ?   :1:  1;
    ?   0   1 (?x) ?   :1:  1;
    *   0   1   x  ?   :1:  1;

    ?   ?   ?   ?  *   :?:  x;

endtable
`endprotect
endprimitive 
// 13 Mar 2002 : Modified such that clrz is dominant than prez, when
//               both the signals are asserted.  In ASIC model
//               prez was dominant.
// 19 Dec 2006 : Sharavathi : changed the timescale for functiononly option to 
//                            1ns/1ps
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
	`timescale	1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module LH100 (  Y );

// Verilog Port Declaration section

   inout  Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

     buf   TI_BUF_PRIM0 ( ACC_Y, Y ) ;


`ifdef TI_functiononly
`else

specify


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//v2.0 03-oct-2009 Guruprasad : Added the behaviourial description.
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module LSR20 (RZ , SZ, Q, QZ ) ;

// Verilog Port Declaration section

   input RZ;
   input SZ;
   output Q;
   output QZ;

`ifdef TETRAMAX

  _DLAT L1 (!SZ,!RZ,1'b0,1'b0,QINT);
  _INV  I1 (QINT, QZINT);
  _OR   O1 (SZ,RZ, SZ_OR_RZ);
  _AND  A1 (SZ_OR_RZ, QINT, Q);
  _AND  A2 (SZ_OR_RZ, QZINT, QZ);

`else


`ifdef TI_verilog    
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     parameter Xon = 1;
     wire GVCnotifier;

//  Verilog Notifier declaration section

    reg GVCnotifier_zd ;

// Xon controlability

   and TI_GVCnotifier (GVCnotifier, Xon, GVCnotifier_zd);

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_SZ_SZ ,  GVC_RZ_RZ  ; 

         srudp   TI_SR_UDP0 ( BFONET1, GVC_SZ_SZ, GVC_RZ_RZ, GVCnotifier ) ;
        srudpz   TI_SRZ_UDP0 ( BFONET2, GVC_SZ_SZ, GVC_RZ_RZ, GVCnotifier ) ;


`else

         srudp   TI_SR_UDP1 ( BFONET1, SZ, RZ, GVCnotifier ) ;
        srudpz   TI_SRZ_UDP1 ( BFONET2, SZ, RZ, GVCnotifier ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          buf #1 TI_BUF_PRIM1 ( QZ, BFONET2 ) ;


`else

          buf  TI_BUF_PRIM2 ( Q, BFONET1 ) ;
          buf  TI_BUF_PRIM3 ( QZ, BFONET2 ) ;

`endif

`ifdef TI_verilog

           not TI_NOT_1 ( INV_RZ, GVC_RZ_RZ );
           or  TI_OR_1 ( COND_SZ, INV_RZ, Q );

`endif


`ifdef TI_functiononly


specify
    $recovery(posedge SZ ,posedge RZ ,1 , GVCnotifier_zd );
endspecify

`else

`ifdef TI_verilog

    wire TCHKON_AND_Q;

    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_COND_SZ;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_COND_SZ (NOT_TCHKON_OR_COND_SZ, COND_SZ, TCHKON_INV);

`endif


specify

      (SZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (SZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (RZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (RZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge SZ &&& (TCHKON_NET != 0) , posedge RZ,  5.0: 5.0: 5.0,  5.0: 5.0: 5.0, GVCnotifier_zd ,,, GVC_SZ_SZ, GVC_RZ_RZ ); 
   $setuphold(posedge RZ &&& (TCHKON_NET != 0) , posedge SZ,  5.0: 5.0: 5.0,  5.0: 5.0: 5.0, GVCnotifier_zd ,,, GVC_RZ_RZ, GVC_SZ_SZ ); 
   $width(negedge RZ &&& TCHKON_AND_Q == 1  ,5.0 : 5.0 : 5.0 , 0 , GVCnotifier_zd) ; 
   $width(negedge SZ &&& NOT_TCHKON_OR_COND_SZ == 0  ,5.0 : 5.0 : 5.0 , 0 , GVCnotifier_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

`endif // ifdef TETRAMAX
endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 09-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module LSR21 (R , S, Q, QZ ) ;

// Verilog Port Declaration section

   input R;
   input S;
   output Q;
   output QZ;

`ifdef TETRAMAX

  _DLAT L1 (S,R,1'b0,1'b0,QINT);
  _INV  I1 (QINT, QZINT);
  _AND   A1 (S,R, S_OR_R);
  _OR  O1 (S_OR_R, QINT, Q);
  _OR  O2 (S_OR_R, QZINT, QZ);

`else


`ifdef TI_verilog    
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     parameter Xon = 1;
     wire GVCnotifier;

//  Verilog Notifier declaration section

    reg GVCnotifier_zd ;

// Xon controlability

   and TI_GVCnotifier (GVCnotifier, Xon, GVCnotifier_zd);

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_S_S ,  GVC_R_R  ; 
	 
         srudp_21   TI_SR_UDP0 ( BFONET1, GVC_S_S, GVC_R_R, GVCnotifier ) ;
        srudpz_21   TI_SRZ_UDP0 ( BFONET2, GVC_S_S, GVC_R_R, GVCnotifier ) ;


`else

         srudp_21   TI_SR_UDP1 ( BFONET1, S, R, GVCnotifier ) ;
        srudpz_21   TI_SRZ_UDP1 ( BFONET2, S, R, GVCnotifier ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          buf #1 TI_BUF_PRIM1 ( QZ, BFONET2 ) ;


`else

          buf  TI_BUF_PRIM2 ( Q, BFONET1 ) ;
          buf  TI_BUF_PRIM3 ( QZ, BFONET2 ) ;

`endif

`ifdef TI_verilog

           not TI_NOT_1 ( INV_S, GVC_S_S );
           and  TI_OR_1 ( COND_R, INV_S, Q );

`endif


`ifdef TI_functiononly


specify
    $recovery(negedge S ,negedge R ,1 , GVCnotifier_zd );
endspecify

`else

`ifdef TI_verilog

    wire TCHKON_AND_Q;
    wire TCHKON_AND_COND_R;

    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_COND_R (TCHKON_AND_COND_R, COND_R, TCHKON_NET);

`endif


specify

      (S *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (S *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (R *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (R *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(negedge S &&& (TCHKON_NET != 0) , negedge R,  5.0: 5.0: 5.0,  5.0: 5.0: 5.0, GVCnotifier_zd ,,, GVC_S_S, GVC_R_R ); 
   $setuphold(negedge R &&& (TCHKON_NET != 0) , negedge S,  5.0: 5.0: 5.0,  5.0: 5.0: 5.0, GVCnotifier_zd ,,, GVC_R_R, GVC_S_S ); 
   $width(posedge R &&& TCHKON_AND_COND_R == 1  ,5.0 : 5.0 : 5.0 , 0 , GVCnotifier_zd) ; 
   $width(posedge S &&& TCHKON_AND_Q == 0  ,5.0 : 5.0 : 5.0 , 0 , GVCnotifier_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

`endif // ifdef TETRAMAX
endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 09-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module MU110F ( A, B, S, Y ) ;

   // Verilog Port Declaration section
        output Y ;
        input A ;
        input B ;
        input S ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        mu1udp #0 TI_MU1UDP_UDP0 ( Y, S, A, B );
        
  `ifdef TI_functiononly

`else
      specify
                ( A *> Y ) = ( 0.0100, 0.0100 ) ;
                ( B *> Y ) = ( 0.0100, 0.0100 ) ;
             if (!A && B)
                ( S *> Y ) = ( 0.0100, 0.0100 ) ;
             if (A && !B)
                ( S *> Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module MU110 ( A, B, S, Y ) ;

   // Verilog Port Declaration section
        output Y ;
        input A ;
        input B ;
        input S ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        mu1udp #0 TI_MU1UDP_UDP0 ( Y, S, A, B );
        
  `ifdef TI_functiononly

`else
      specify
                ( A *> Y ) = ( 0.0100, 0.0100 ) ;
                ( B *> Y ) = ( 0.0100, 0.0100 ) ;
             if (!A && B)
                ( S *> Y ) = ( 0.0100, 0.0100 ) ;
             if (A && !B)
                ( S *> Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module MU111 ( AZ, B, S, Y ) ;

  // Verilog Port Declaration section
        output Y ;
        input AZ ;
        input B ;
        input S ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not TI_NOT_PRIM0 ( A, AZ );
        mu1udp #0 TI_MU1UDP_UDP0  ( Y, S, A, B );
`ifdef TI_functiononly

`else

        specify
                ( AZ *> Y ) = ( 0.0100, 0.0100 ) ;
                ( B *> Y ) = ( 0.0100, 0.0100 ) ;
             if (AZ && B)
                ( S *> Y ) = ( 0.0100, 0.0100 ) ;
             if (!AZ && !B)
                ( S *> Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module MU112 ( A, B, S, YZ ) ;

  // Verilog Port Declaration section
        output YZ ;
        input A ;
        input B ;
        input S ;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
        mu1udp TI_MU1UDP_UDP0 ( Y, S, A, B );
        not #0 TI_NOT_PRIM0 ( YZ, Y );

`ifdef TI_functiononly

`else
        specify
                ( A *> YZ ) = ( 0.0100, 0.0100 ) ;
                ( B *> YZ ) = ( 0.0100, 0.0100 ) ;
             if (!A && B)
                ( S *> YZ ) = ( 0.0100, 0.0100 ) ;
             if (A && !B)
                ( S *> YZ ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module MU120F ( A, B, S, Y ) ;

   // Verilog Port Declaration section
        output Y ;
        input A ;
        input B ;
        input S ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        mu1udp #0 TI_MU1UDP_UDP0 ( Y, S, A, B );
        
  `ifdef TI_functiononly

`else
      specify
                ( A *> Y ) = ( 0.0100, 0.0100 ) ;
                ( B *> Y ) = ( 0.0100, 0.0100 ) ;
             if (!A && B)
                ( S *> Y ) = ( 0.0100, 0.0100 ) ;
             if (A && !B)
                ( S *> Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module MU120 ( A, B, S, Y ) ;

   // Verilog Port Declaration section
        output Y ;
        input A ;
        input B ;
        input S ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        mu1udp #0 TI_MU1UDP_UDP0 ( Y, S, A, B );
        
  `ifdef TI_functiononly

`else
      specify
                ( A *> Y ) = ( 0.0100, 0.0100 ) ;
                ( B *> Y ) = ( 0.0100, 0.0100 ) ;
             if (!A && B)
                ( S *> Y ) = ( 0.0100, 0.0100 ) ;
             if (A && !B)
                ( S *> Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module MU122 ( A, B, S, YZ ) ;

  // Verilog Port Declaration section
        output YZ ;
        input A ;
        input B ;
        input S ;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
        mu1udp TI_MU1UDP_UDP0 ( Y, S, A, B );
        not #0 TI_NOT_PRIM0 ( YZ, Y );

`ifdef TI_functiononly

`else
        specify
                ( A *> YZ ) = ( 0.0100, 0.0100 ) ;
                ( B *> YZ ) = ( 0.0100, 0.0100 ) ;
             if (!A && B)
                ( S *> YZ ) = ( 0.0100, 0.0100 ) ;
             if (A && !B)
                ( S *> YZ ) = ( 0.0100, 0.0100 ) ;
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif



// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module MU140F ( A, B, S, Y ) ;

   // Verilog Port Declaration section
        output Y ;
        input A ;
        input B ;
        input S ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        mu1udp #0 TI_MU1UDP_UDP0 ( Y, S, A, B );
        
  `ifdef TI_functiononly

`else
      specify
                ( A *> Y ) = ( 0.0100, 0.0100 ) ;
                ( B *> Y ) = ( 0.0100, 0.0100 ) ;
             if (!A && B)
                ( S *> Y ) = ( 0.0100, 0.0100 ) ;
             if (A && !B)
                ( S *> Y ) = ( 0.0100, 0.0100 ) ;
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2002 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------


`resetall
`ifdef TI_functiononly
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

primitive mu1udp
`protect
(Q, S, A, B);
output Q; 
input S, A, B;

table
//      S  A  B   Q
        0  0  ?  : 0 ;
        0  1  ?  : 1 ;
        0  x  ?  : x ;
        1  ?  0  : 0 ;
        1  ?  1  : 1 ;
        1  ?  x  : x ;
        x  0  0  : 0 ;
        x  1  1  : 1 ;

endtable
`endprotect
endprimitive
// Revision history:
// ----------------
// v1.2  08-Jun-1999  Changing 10ps to 1ps
// v1.1  17-Mar-1999 24 date and time created 99/03/17 17
// 19 Dec 2006 : Sharavathi : changed the timescale for functiononly option to 
//                            1ns/1ps 
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module MU210 ( A, B, C, D, S1, S2, Y ) ;

   // Verilog Port Declaration section
        output Y ;
        input A ;
        input B ;
        input C ;
        input D ;
        input S1 ;
        input S2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        mu2udp #0 TI_MU2UDP_UDP0( Y, S1, S2, A, B, C, D );
  `ifdef TI_functiononly

`else

        specify
             if ( !A && B && !C && !D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && C && !D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && B && C && !D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && C && !D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && !B && C && !D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && !B && !C && D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && !C && D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && B && !C && D && S2  )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && !C && D  && S2)
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && !C && D  && !S2)
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && !C && !D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && C && !D && !S2)
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && C && D && !S2)
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && C && !D && !S2)
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && C && D && !S2)
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && !C && D && !S2)
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && !C && !D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && B && !C && !D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && B && C && !D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && C && !D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && B && !C && D && !S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && B && !C && !D && !S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && !C && !D && !S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
	     if ( !A && !B && !C && D && S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );  
             if (  A && !B && !C && D && !S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && !C && D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A&& !B && C && D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && C && D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && !B && C && D  && !S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && !B && C && !D  && !S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && C && !D  && !S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && C && D  && !S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if (B && !C && !D )
                  ( A *>  Y) = ( 0.0100, 0.0100 );
             if (!B && C && D )
                  ( A *>  Y) = ( 0.0100, 0.0100 );
             if (!B && !C && D )
                  ( A *>  Y) = ( 0.0100, 0.0100 );
             if (!B && !C && !D )
                  ( A *>  Y) = ( 0.0100, 0.0100 );
             if (!B && C && !D )
                  ( A *>  Y) = ( 0.0100, 0.0100 );
             if (B && C && !D )
                  ( A *>  Y) = ( 0.0100, 0.0100 );
             if (B && C && D )
                  ( A *>  Y) = ( 0.0100, 0.0100 );
             if (B && !C && D )
                  ( A *>  Y) = ( 0.0100, 0.0100 );
             if (A && !C && D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (!A && !C && D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (!A && C && D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (!A && C && !D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (!A && !C && !D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (A && !C && !D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (A && C && !D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (A && C && D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (!A && B && !D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (!A && !B && !D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (!A && !B && D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (!A && B && D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (A && B && D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (A && B && !D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (A && !B && !D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (A && !B && D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (!A && B && !C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (A && B && !C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (A && !B && !C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (A && !B && C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (A && B && C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (!A && B && C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (!A && !B && C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (!A && !B && !C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module MU211 ( AZ, B, C, D, S1, S2, Y ) ;

    // Verilog Port Declaration section
        output Y ;
        input AZ ;
        input B ;
        input C ;
        input D ;
        input S1 ;
        input S2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not TI_NOT_PRIM0 ( A, AZ );
        mu2udp #0 TI_MU2UDP_UDP0( Y, S1, S2, A, B, C, D );

 `ifdef TI_functiononly

`else
       specify
             if ( AZ && B && !C && !D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && !B && C && !D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && B && C && !D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && B && C && !D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && !B && C && !D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && !B && !C && D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && B && !C && D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && B && !C && D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && !B && !C && D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && !B && !C && D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && !B && !C && !D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && !B && C && !D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && !B && C && D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && B && C && !D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && B && C && D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && B && !C && D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && B && !C && !D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && B && !C && !D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && B && C && !D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && B && C && !D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && B && !C && D && !S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && B && !C && !D && !S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && !B && !C && !D && !S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && !B && !C && D && !S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && !B && !C && D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && !B && !C && D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && !B && C && D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && !B && C && D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && !B && C && D && !S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && !B && C && !D && !S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && B && C && !D && !S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && B && C && D && !S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if (B && !C && !D )
                  ( AZ *>  Y) = ( 0.0100, 0.0100 );
             if (!B && C && D )
                  ( AZ *>  Y) = ( 0.0100, 0.0100 );
             if (!B && !C && D )
                  ( AZ *>  Y) = ( 0.0100, 0.0100 );
             if (!B && !C && !D )
                  ( AZ *>  Y) = ( 0.0100, 0.0100 );
             if (!B && C && !D )
                  ( AZ *>  Y) = ( 0.0100, 0.0100 );
             if (B && C && !D )
                  ( AZ *>  Y) = ( 0.0100, 0.0100 );
             if (B && C && D )
                  ( AZ *>  Y) = ( 0.0100, 0.0100 );
             if (B && !C && D )
                  ( AZ *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && !C && D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && !C && D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && C && D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && C && !D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && !C && !D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && !C && !D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && C && !D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && C && D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && B && !D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && !B && !D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && !B && D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && B && D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && B && D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && B && !D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && !B && !D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && !B && D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && B && !C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && B && !C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && !B && !C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && !B && C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && B && C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && B && C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && !B && C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && !B && !C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module MU212 ( AZ, BZ, C, D, S1, S2, Y ) ;

    // Verilog Port Declaration section
        output Y ;
        input AZ ;
        input BZ ;
        input C ;
        input D ;
        input S1 ;
        input S2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not TI_NOT_PRIM0 ( A, AZ );
        not TI_NOT_PRIM1 ( B, BZ );
        mu2udp #0  TI_MU2UDP_UDP0 ( Y, S1, S2, A, B, C, D );
`ifdef TI_functiononly

`else


        specify
             if ( AZ && !BZ && !C && !D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && BZ && C && !D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && !BZ && C && !D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && !BZ && C && !D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && BZ && C && !D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && BZ && !C && D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && !BZ && !C && D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && !BZ && !C && D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && BZ && !C && D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && BZ && !C && D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && BZ && !C && !D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && BZ && C && !D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && BZ && C && D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && !BZ && C && !D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && !BZ && C && D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && !BZ && !C && D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && !BZ && !C && !D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && !BZ && !C && !D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && !BZ && C && !D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && !BZ && C && !D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && !BZ && !C && D && !S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && !BZ && !C && !D && !S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && BZ && !C && !D && !S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && BZ && !C && D && !S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && BZ && !C && D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && BZ && !C && D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && BZ && C && D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !AZ && BZ && C && D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && BZ && C && D && !S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && BZ && C && !D && !S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && !BZ && C && !D && !S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( AZ && !BZ && C && D && !S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if (!BZ && !C && !D )
                  ( AZ *>  Y) = ( 0.0100, 0.0100 );
             if (BZ && C && D )
                  ( AZ *>  Y) = ( 0.0100, 0.0100 );
             if (BZ && !C && D )
                  ( AZ *>  Y) = ( 0.0100, 0.0100 );
             if (BZ && !C && !D )
                  ( AZ *>  Y) = ( 0.0100, 0.0100 );
             if (BZ && C && !D )
                  ( AZ *>  Y) = ( 0.0100, 0.0100 );
             if (!BZ && C && !D )
                  ( AZ *>  Y) = ( 0.0100, 0.0100 );
             if (!BZ && C && D )
                  ( AZ *>  Y) = ( 0.0100, 0.0100 );
             if (!BZ && !C && D )
                  ( AZ *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && !C && D )
                  ( BZ *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && !C && D )
                  ( BZ *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && C && D )
                  ( BZ *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && C && !D )
                  ( BZ *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && !C && !D )
                  ( BZ *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && !C && !D )
                  ( BZ *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && C && !D )
                  ( BZ *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && C && D )
                  ( BZ *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && !BZ && !D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && BZ && !D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && BZ && D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && !BZ && D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && !BZ && D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && !BZ && !D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && BZ && !D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && BZ && D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && !BZ && !C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && !BZ && !C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && BZ && !C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && BZ && C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (!AZ && !BZ && C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && !BZ && C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && BZ && C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (AZ && BZ && !C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
        endspecify


`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module MU214 ( A, B, C, D, S1, S2, YZ ) ;

   // Verilog Port Declaration section
        output YZ ;
        input A ;
        input B ;
        input C ;
        input D ;
        input S1 ;
        input S2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        mu2udp TI_MU2UDP_UDP0 ( Y, S1, S2, A, B, C, D );
        not #0 TI_NOT_PRIM0 ( YZ, Y );

     `ifdef TI_functiononly

`else
     specify
             if ( !A && B && !C && !D && !S2 )
                  ( S1 *>  YZ) = ( 0.0100, 0.0100 );
             if ( A && !B && C && !D && S2 )
                  ( S1 *>  YZ) = ( 0.0100, 0.0100 );
             if ( A && B && C && !D && S2 )
                  ( S1 *>  YZ) = ( 0.0100, 0.0100 );
             if ( !A && B && C && !D && S2 )
                  ( S1 *>  YZ) = ( 0.0100, 0.0100 );
             if ( !A && !B && C && !D && S2 )
                  ( S1 *>  YZ) = ( 0.0100, 0.0100 );
             if ( !A && !B && !C && D && S2 )
                  ( S1 *>  YZ) = ( 0.0100, 0.0100 );
             if ( !A && B && !C && D && S2 )
                  ( S1 *>  YZ) = ( 0.0100, 0.0100 );
             if ( A && B && !C && D && S2 )
                  ( S1 *>  YZ) = ( 0.0100, 0.0100 );
             if ( A && !B && !C && D && S2 )
                  ( S1 *>  YZ) = ( 0.0100, 0.0100 );
             if ( A && !B && !C && D && !S2 )
                  ( S1 *>  YZ) = ( 0.0100, 0.0100 );
             if ( A && !B && !C && !D && !S2 )
                  ( S1 *>  YZ) = ( 0.0100, 0.0100 );
             if ( A && !B && C && !D && !S2 )
                  ( S1 *>  YZ) = ( 0.0100, 0.0100 );
             if ( A && !B && C && D && !S2 )
                  ( S1 *>  YZ) = ( 0.0100, 0.0100 );
             if ( !A && B && C && !D && !S2 )
                  ( S1 *>  YZ) = ( 0.0100, 0.0100 );
             if ( !A && B && C && D && !S2 )
                  ( S1 *>  YZ) = ( 0.0100, 0.0100 );
             if ( !A && B && !C && D && !S2 )
                  ( S1 *>  YZ) = ( 0.0100, 0.0100 );
             if ( !A && B && !C && !D && S1 )
                  ( S2 *>  YZ) = ( 0.0100, 0.0100 );
             if ( A && B && !C && !D && S1 )
                  ( S2 *>  YZ) = ( 0.0100, 0.0100 );
             if ( A && B && C && !D && S1 )
                  ( S2 *>  YZ) = ( 0.0100, 0.0100 );
             if ( !A && B && C && !D && S1 )
                  ( S2 *>  YZ) = ( 0.0100, 0.0100 );
             if ( A && B && !C && D && !S1 )
                  ( S2 *>  YZ) = ( 0.0100, 0.0100 );
             if ( A && B && !C && !D && !S1 )
                  ( S2 *>  YZ) = ( 0.0100, 0.0100 );
             if ( A && !B && !C && !D && !S1 )
                  ( S2 *>  YZ) = ( 0.0100, 0.0100 );
             if ( A && !B && !C && D && !S1 )
                  ( S2 *>  YZ) = ( 0.0100, 0.0100 );
             if ( A && !B && !C && D && S1 )
                  ( S2 *>  YZ) = ( 0.0100, 0.0100 );
             if ( !A && !B && !C && D && S1 )
                  ( S2 *>  YZ) = ( 0.0100, 0.0100 );
             if ( !A && !B && C && D && S1 )
                  ( S2 *>  YZ) = ( 0.0100, 0.0100 );
             if ( A && !B && C && D && S1 )
                  ( S2 *>  YZ) = ( 0.0100, 0.0100 );
             if ( !A && !B && C && D && !S1 )
                  ( S2 *>  YZ) = ( 0.0100, 0.0100 );
             if ( !A && !B && C && !D && !S1 )
                  ( S2 *>  YZ) = ( 0.0100, 0.0100 );
             if ( !A && B && C && !D && !S1 )
                  ( S2 *>  YZ) = ( 0.0100, 0.0100 );
             if ( !A && B && C && D && !S1 )
                  ( S2 *>  YZ) = ( 0.0100, 0.0100 );
             if (B && !C && !D )
                  ( A *>  YZ) = ( 0.0100, 0.0100 );
             if (!B && C && D )
                  ( A *>  YZ) = ( 0.0100, 0.0100 );
             if (!B && !C && D )
                  ( A *>  YZ) = ( 0.0100, 0.0100 );
             if (!B && !C && !D )
                  ( A *>  YZ) = ( 0.0100, 0.0100 );
             if (!B && C && !D )
                  ( A *>  YZ) = ( 0.0100, 0.0100 );
             if (B && C && !D )
                  ( A *>  YZ) = ( 0.0100, 0.0100 );
             if (B && C && D )
                  ( A *>  YZ) = ( 0.0100, 0.0100 );
             if (B && !C && D )
                  ( A *>  YZ) = ( 0.0100, 0.0100 );
             if (A && !C && D )
                  ( B *>  YZ) = ( 0.0100, 0.0100 );
             if (!A && !C && D )
                  ( B *>  YZ) = ( 0.0100, 0.0100 );
             if (!A && C && D )
                  ( B *>  YZ) = ( 0.0100, 0.0100 );
             if (!A && C && !D )
                  ( B *>  YZ) = ( 0.0100, 0.0100 );
             if (!A && !C && !D )
                  ( B *>  YZ) = ( 0.0100, 0.0100 );
             if (A && !C && !D )
                  ( B *>  YZ) = ( 0.0100, 0.0100 );
             if (A && C && !D )
                  ( B *>  YZ) = ( 0.0100, 0.0100 );
             if (A && C && D )
                  ( B *>  YZ) = ( 0.0100, 0.0100 );
             if (!A && B && !D )
                  ( C *>  YZ) = ( 0.0100, 0.0100 );
             if (!A && !B && !D )
                  ( C *>  YZ) = ( 0.0100, 0.0100 );
             if (!A && !B && D )
                  ( C *>  YZ) = ( 0.0100, 0.0100 );
             if (!A && B && D )
                  ( C *>  YZ) = ( 0.0100, 0.0100 );
             if (A && B && D )
                  ( C *>  YZ) = ( 0.0100, 0.0100 );
             if (A && B && !D )
                  ( C *>  YZ) = ( 0.0100, 0.0100 );
             if (A && !B && !D )
                  ( C *>  YZ) = ( 0.0100, 0.0100 );
             if (A && !B && D )
                  ( C *>  YZ) = ( 0.0100, 0.0100 );
             if (!A && B && !C )
                  ( D *>  YZ) = ( 0.0100, 0.0100 );
             if (A && B && !C )
                  ( D *>  YZ) = ( 0.0100, 0.0100 );
             if (A && !B && !C )
                  ( D *>  YZ) = ( 0.0100, 0.0100 );
             if (A && !B && C )
                  ( D *>  YZ) = ( 0.0100, 0.0100 );
             if (A && B && C )
                  ( D *>  YZ) = ( 0.0100, 0.0100 );
             if (!A && B && C )
                  ( D *>  YZ) = ( 0.0100, 0.0100 );
             if (!A && !B && C )
                  ( D *>  YZ) = ( 0.0100, 0.0100 );
             if (!A && !B && !C )
                  ( D *>  YZ) = ( 0.0100, 0.0100 );
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module MU220 ( A, B, C, D, S1, S2, Y ) ;

   // Verilog Port Declaration section
        output Y ;
        input A ;
        input B ;
        input C ;
        input D ;
        input S1 ;
        input S2 ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        mu2udp #0 TI_MU2UDP_UDP0( Y, S1, S2, A, B, C, D );
  `ifdef TI_functiononly

`else

        specify
             if ( !A && B && !C && !D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && C && !D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && B && C && !D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && C && !D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && !B && C && !D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && !B && !C && D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && !C && D && S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && B && !C && D && S2  )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && !C && D  && S2)
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && !C && D  && !S2)
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && !C && !D && !S2 )
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && C && !D && !S2)
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && C && D && !S2)
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && C && !D && !S2)
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && C && D && !S2)
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && !C && D && !S2)
                  ( S1 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && !C && !D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && B && !C && !D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && B && C && !D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && C && !D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && B && !C && D && !S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && B && !C && !D && !S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && !C && !D && !S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
	     if ( !A && !B && !C && D && S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );  
             if (  A && !B && !C && D && !S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && !C && D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A&& !B && C && D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( A && !B && C && D && S1 )
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && !B && C && D  && !S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && !B && C && !D  && !S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && C && !D  && !S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if ( !A && B && C && D  && !S1)
                  ( S2 *>  Y) = ( 0.0100, 0.0100 );
             if (B && !C && !D )
                  ( A *>  Y) = ( 0.0100, 0.0100 );
             if (!B && C && D )
                  ( A *>  Y) = ( 0.0100, 0.0100 );
             if (!B && !C && D )
                  ( A *>  Y) = ( 0.0100, 0.0100 );
             if (!B && !C && !D )
                  ( A *>  Y) = ( 0.0100, 0.0100 );
             if (!B && C && !D )
                  ( A *>  Y) = ( 0.0100, 0.0100 );
             if (B && C && !D )
                  ( A *>  Y) = ( 0.0100, 0.0100 );
             if (B && C && D )
                  ( A *>  Y) = ( 0.0100, 0.0100 );
             if (B && !C && D )
                  ( A *>  Y) = ( 0.0100, 0.0100 );
             if (A && !C && D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (!A && !C && D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (!A && C && D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (!A && C && !D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (!A && !C && !D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (A && !C && !D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (A && C && !D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (A && C && D )
                  ( B *>  Y) = ( 0.0100, 0.0100 );
             if (!A && B && !D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (!A && !B && !D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (!A && !B && D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (!A && B && D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (A && B && D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (A && B && !D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (A && !B && !D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (A && !B && D )
                  ( C *>  Y) = ( 0.0100, 0.0100 );
             if (!A && B && !C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (A && B && !C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (A && !B && !C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (A && !B && C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (A && B && C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (!A && B && C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (!A && !B && C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
             if (!A && !B && !C )
                  ( D *>  Y) = ( 0.0100, 0.0100 );
        endspecify

`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
// mu2udp.v - verilog model

`resetall
`ifdef TI_functiononly
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

primitive mu2udp
`protect
(y, s1, s2, a, b, c, d);
    output y;
//    reg y;    
    input s1, s2, a, b, c, d;
    
    table   
//      s1  s2  a   b   c   d    y
        0   0   1   ?   ?   ?  : 1  ;
        0   0   0   ?   ?   ?  : 0  ;
        0   0   x   ?   ?   ?  : x  ;
        1   0   ?   1   ?   ?  : 1  ;
        1   0   ?   0   ?   ?  : 0  ;
        1   0   ?   x   ?   ?  : x  ;
        0   1   ?   ?   1   ?  : 1  ;
        0   1   ?   ?   0   ?  : 0  ;
        0   1   ?   ?   x   ?  : x  ;
        1   1   ?   ?   ?   1  : 1  ;
        1   1   ?   ?   ?   0  : 0  ;
        1   1   ?   ?   ?   x  : x  ;
        x   0   1   1   ?   ?  : 1  ;
        x   0   0   0   ?   ?  : 0  ;
        x   1   ?   ?   1   1  : 1  ;
        x   1   ?   ?   0   0  : 0  ;
        0   x   1   ?   1   ?  : 1  ;
        0   x   0   ?   0   ?  : 0  ;
        1   x   ?   1   ?   1  : 1  ;
        1   x   ?   0   ?   0  : 0  ;
        x   x   0   0   0   0  : 0  ;
        x   x   1   1   1   1  : 1  ;

    endtable

`endprotect

endprimitive 

// 19 Dec 2006 : Sharavathi : changed the timescale for functiononly option to 
//                            1ns/1ps

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
// 21-Jan-2010 Mazhar. Updated to add timescale in TI-functiononly with 
//             if else statement and add resetall statement
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA210F (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA210 (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NA211F (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nand #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NA211 (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nand #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA220F (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA220 (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NA221F (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nand #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NA221 (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nand #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA240F (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA240 (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NA241F (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nand #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NA241 (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nand #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA260F (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NA261F (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nand #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA280F (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA310F (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA310 (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NA311F (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nand #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NA311 (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nand #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA320F (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA320 (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NA321F (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nand #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NA321 (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nand #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA340F (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA340 (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NA341F (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nand #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NA341 (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nand #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA360F (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NA361F (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nand #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA380F (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA410F (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA410 (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module NA411 ( AZ, B, C, D, Y ) ;

 // Verilog Port Declaration section
        output Y ;
        input AZ ;
        input B ;
        input C ;
        input D ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
      not TI_NOT_PRIM0 ( A, AZ );
      nand #0 TI_NAND_PRIM0 ( Y, A, B, C, D ) ;
`ifdef TI_functiononly
`else

        specify
                ( AZ => Y ) = ( 0.0100, 0.0100 ) ;
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
                ( C => Y ) = ( 0.0100, 0.0100 ) ;
                ( D => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA420F (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA420 (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module NA421 ( AZ, B, C, D, Y ) ;

 // Verilog Port Declaration section
        output Y ;
        input AZ ;
        input B ;
        input C ;
        input D ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
      not TI_NOT_PRIM0 ( A, AZ );
      nand #0 TI_NAND_PRIM0 ( Y, A, B, C, D ) ;
`ifdef TI_functiononly
`else

        specify
                ( AZ => Y ) = ( 0.0100, 0.0100 ) ;
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
                ( C => Y ) = ( 0.0100, 0.0100 ) ;
                ( D => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA440F (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA440 (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module NA441 ( AZ, B, C, D, Y ) ;

 // Verilog Port Declaration section
        output Y ;
        input AZ ;
        input B ;
        input C ;
        input D ;

  `ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
      not TI_NOT_PRIM0 ( A, AZ );
      nand #0 TI_NAND_PRIM0 ( Y, A, B, C, D ) ;
`ifdef TI_functiononly
`else

        specify
                ( AZ => Y ) = ( 0.0100, 0.0100 ) ;
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
                ( C => Y ) = ( 0.0100, 0.0100 ) ;
                ( D => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NA460F (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nand #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO210F (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO210 (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NO211F (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nor #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NO211 (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nor #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO220F (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO220 (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NO221F (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nor #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NO221 (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nor #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO240F (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO240 (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NO241F (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nor #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NO241 (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nor #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO260F (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NO261F (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nor #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO310F (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO310 (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NO311F (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nor #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NO311 (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nor #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO320F (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO320 (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NO321F (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nor #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NO321 (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nor #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO340F (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO340 (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NO341F (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nor #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NO341 (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nor #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO360F (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module  NO361F (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           nor #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO410 (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module NO411 ( AZ, B, C, D, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input AZ ;
        input B ;
        input C ;
        input D ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not TI_NOT_PRIM0 ( A, AZ );
        nor #0 TI_NOR_PRIM0 ( Y, A, B, C, D ) ;

 `ifdef TI_functiononly
`else
       specify
                ( AZ => Y ) = ( 0.0100, 0.0100 ) ;
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
                ( C => Y ) = ( 0.0100, 0.0100 ) ;
                ( D => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO420 (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module NO421 ( AZ, B, C, D, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input AZ ;
        input B ;
        input C ;
        input D ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not TI_NOT_PRIM0 ( A, AZ );
        nor #0 TI_NOR_PRIM0 ( Y, A, B, C, D ) ;

 `ifdef TI_functiononly
`else
       specify
                ( AZ => Y ) = ( 0.0100, 0.0100 ) ;
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
                ( C => Y ) = ( 0.0100, 0.0100 ) ;
                ( D => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module  NO440 (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           nor #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module NO441 ( AZ, B, C, D, Y ) ;

// Verilog Port Declaration section
        output Y ;
        input AZ ;
        input B ;
        input C ;
        input D ;
`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

        not TI_NOT_PRIM0 ( A, AZ );
        nor #0 TI_NOR_PRIM0 ( Y, A, B, C, D ) ;

 `ifdef TI_functiononly
`else
       specify
                ( AZ => Y ) = ( 0.0100, 0.0100 ) ;
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
                ( C => Y ) = ( 0.0100, 0.0100 ) ;
                ( D => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module OR210 (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           or #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module OR211 (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           or #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module OR220 (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           or #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module OR221 (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           or #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module OR240 (  A , B , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           or #0 TI_AND_PRIM0 ( Y , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module OR241 (AZ , B, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           or #0 TI_AND_PRIM0 ( Y, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module OR310 (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           or #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module OR311 (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           or #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module OR320 (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           or #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module OR321 (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           or #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module OR340 (  A , B , C , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           or #0 TI_AND_PRIM0 ( Y , C , A , B ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module OR341 (AZ , B, C, Y ) ;

// Verilog Port Declaration section

   input AZ;
   input B;
   input C;
   output Y;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

 
           not   TI_NOT_PRIM0 ( IINVnet1, AZ ) ;
           or #0 TI_AND_PRIM0 ( Y, C, IINVnet1, B ) ;


`ifdef TI_functiononly

`else


specify

    (AZ -=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (B +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);
    (C +=> Y) = (0.010000:0.010000:0.010000 , 0.010000:0.010000:0.010000);


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module OR410 (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           or #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module OR411 ( AZ, B, C, D, Y ) ;

   // Verilog Port Declaration section
     output Y ;
        input AZ ;
        input B ;
        input C ;
        input D ;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
        not TI_NOT_PRIM0  ( A, AZ );
           or #0 TI_OR_PRIM0 ( Y, A, B, C, D ) ;

 `ifdef TI_functiononly
`else
       specify
                ( AZ => Y ) = ( 0.0100, 0.0100 ) ;
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
                ( C => Y ) = ( 0.0100, 0.0100 ) ;
                ( D => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module OR420 (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           or #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module OR421 ( AZ, B, C, D, Y ) ;

   // Verilog Port Declaration section
     output Y ;
        input AZ ;
        input B ;
        input C ;
        input D ;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
        not TI_NOT_PRIM0  ( A, AZ );
           or #0 TI_OR_PRIM0 ( Y, A, B, C, D ) ;

 `ifdef TI_functiononly
`else
       specify
                ( AZ => Y ) = ( 0.0100, 0.0100 ) ;
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
                ( C => Y ) = ( 0.0100, 0.0100 ) ;
                ( D => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module OR440 (  A , B , C , D , Y );

// Verilog Port Declaration section

   input  A;
   input  B;
   input  C;
   input  D;
   output Y;


`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)


           or #0 TI_AND_PRIM0 ( Y , A , B , C , D ) ;

`ifdef TI_functiononly
`else

specify

    (A +=> Y)  = 0.01 ;
    (B +=> Y)  = 0.01 ;
    (C +=> Y)  = 0.01 ;
    (D +=> Y)  = 0.01 ;

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif
// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine


`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module OR441 ( AZ, B, C, D, Y ) ;

   // Verilog Port Declaration section
     output Y ;
        input AZ ;
        input B ;
        input C ;
        input D ;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)
        not TI_NOT_PRIM0  ( A, AZ );
           or #0 TI_OR_PRIM0 ( Y, A, B, C, D ) ;

 `ifdef TI_functiononly
`else
       specify
                ( AZ => Y ) = ( 0.0100, 0.0100 ) ;
                ( B => Y ) = ( 0.0100, 0.0100 ) ;
                ( C => Y ) = ( 0.0100, 0.0100 ) ;
                ( D => Y ) = ( 0.0100, 0.0100 ) ;
        endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module SDB20 (CLK , CLRZ, D, PREZ, S, SD, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input PREZ;
   input S;
   input SD;
   output Q;
   output QZ;

`ifdef TETRAMAX
   _INV I1  ( CLRZ,CLR);
   _INV I2  ( PREZ,PRE);
   _NAND N1 ( CLR,PRE,CLR_PRE);
   _MUX M2  ( S, D, SD, DINT );
   _DFF FF1 ( !PREZ, !CLRZ, CLK, DINT, QINT);
   _INV I3  ( QINT,QZINT);
   _AND A1  ( CLRZ,QINT,Q1);
   _AND A2  ( PRE,CLR_PRE,Q2);
   _AND A3  ( QZINT,PREZ, Q3);
   _AND A4  ( CLR, CLR_PRE, Q4);
   _OR  O1  ( Q1,Q2,Q);
   _OR  O2  ( Q3,Q4,QZ);
`else
 


`ifdef TI_verilog    
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     parameter Xon = 1;
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_CLRZ_CLRZ  ,  GVC_PREZ_PREZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
        dlaudp   TI_DLA_UDP0 ( FNET4, DIN, IINVnet1, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP1 ( BFONET1, FNET4, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP0 ( BFONET2, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, BFONET1 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
        dlaudp   TI_DLA_UDP2 ( FNET4, DIN, IINVnet1, CLRZ, PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP3 ( BFONET1, FNET4, CLK, CLRZ, PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP1 ( BFONET2, CLRZ, PREZ, BFONET1 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          buf #1 TI_BUF_PRIM1 ( QZ, BFONET2 ) ;


`else

          buf  TI_BUF_PRIM2 ( Q, BFONET1 ) ;
          buf  TI_BUF_PRIM3 ( QZ, BFONET2 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ , 1'b0 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND4 ( GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ , 1'b1 , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND5 ( GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND6 ( GVC_Q_NOT0_PREZ_NOT0_ , Q , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND7 ( GVC_Q_NOT1_CLRZ_NOT0_ , Q , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly


specify
    $recovery(posedge PREZ ,posedge CLRZ ,1 , GVCnotifier2_zd );
endspecify

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_;

    and TI_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_, GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_, GVC_Q_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_, GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_, GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ (TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_, GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_, GVC_Q_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_, GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ (TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_, GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_, TCHKON_NET);

`endif


specify
      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ != 0  , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $setuphold(posedge PREZ &&& (TCHKON_NET != 0) , posedge CLRZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_PREZ_PREZ, GVC_CLRZ_CLRZ ); 
   $setuphold(posedge CLRZ &&& (TCHKON_NET != 0) , posedge PREZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ  &&& TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge PREZ  &&& TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

`endif // ifdef TETRAMAX
endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 09-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module SDB23 (CLK , CLRZ, D, PREZ, S, SD, Q ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input PREZ;
   input S;
   input SD;
   output Q;

`ifdef TETRAMAX
   _INV I1  ( CLRZ,CLR);
   _INV I2  ( PREZ,PRE);
   _NAND N1 ( CLR,PRE,CLR_PRE);
   _MUX M2  ( S, D, SD, DINT );
   _DFF FF1 ( !PREZ, !CLRZ, CLK, DINT, QINT);
   _INV I3  ( QINT,QZINT);
   _AND A1  ( CLRZ,QINT,Q1);
   _AND A2  ( PRE,CLR_PRE,Q2);
   _AND A3  ( QZINT,PREZ, Q3);
   _AND A4  ( CLR, CLR_PRE, Q4);
   _OR  O1  ( Q1,Q2,Q);
`else
 


`ifdef TI_verilog    
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     parameter Xon = 1;
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_CLRZ_CLRZ  ,  GVC_PREZ_PREZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
        dlaudp   TI_DLA_UDP0 ( FNET4, DIN, IINVnet1, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP1 ( BFONET1, FNET4, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP0 ( BFONET2, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, BFONET1 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
        dlaudp   TI_DLA_UDP2 ( FNET4, DIN, IINVnet1, CLRZ, PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP3 ( BFONET1, FNET4, CLK, CLRZ, PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP1 ( BFONET2, CLRZ, PREZ, BFONET1 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          buf  TI_BUF_PRIM1 ( QZ, BFONET2 ) ;


`else

          buf  TI_BUF_PRIM2 ( Q, BFONET1 ) ;
          buf  TI_BUF_PRIM3 ( QZ, BFONET2 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ , 1'b0 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND4 ( GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ , 1'b1 , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND5 ( GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND6 ( GVC_Q_NOT0_PREZ_NOT0_ , Q , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND7 ( GVC_Q_NOT1_CLRZ_NOT0_ , Q , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly


specify
    $recovery(posedge PREZ ,posedge CLRZ ,1 , GVCnotifier2_zd );
endspecify

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_;

    and TI_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_, GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_, GVC_Q_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_, GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_, GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ (TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_, GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_, GVC_Q_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_, GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ (TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_, GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_, TCHKON_NET);

`endif


specify
      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ != 0  , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $setuphold(posedge PREZ &&& (TCHKON_NET != 0) , posedge CLRZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_PREZ_PREZ, GVC_CLRZ_CLRZ ); 
   $setuphold(posedge CLRZ &&& (TCHKON_NET != 0) , posedge PREZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ  &&& TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge PREZ  &&& TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

`endif // ifdef TETRAMAX
endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 09-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module SDB24 (CLK , CLRZ, D, PREZ, S, SD,  QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input PREZ;
   input S;
   input SD;
   output QZ;

`ifdef TETRAMAX
   _INV I1  ( CLRZ,CLR);
   _INV I2  ( PREZ,PRE);
   _NAND N1 ( CLR,PRE,CLR_PRE);
   _MUX M2  ( S, D, SD, DINT );
   _DFF FF1 ( !PREZ, !CLRZ, CLK, DINT, QINT);
   _INV I3  ( QINT,QZINT);
   _AND A1  ( CLRZ,QINT,Q1);
   _AND A2  ( PRE,CLR_PRE,Q2);
   _AND A3  ( QZINT,PREZ, Q3);
   _AND A4  ( CLR, CLR_PRE, Q4);
   _OR  O2  ( Q3,Q4,QZ);
`else
 


`ifdef TI_verilog    
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     parameter Xon = 1;
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_CLRZ_CLRZ  ,  GVC_PREZ_PREZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
        dlaudp   TI_DLA_UDP0 ( FNET4, DIN, IINVnet1, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP1 ( BFONET1, FNET4, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP0 ( BFONET2, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, BFONET1 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
        dlaudp   TI_DLA_UDP2 ( FNET4, DIN, IINVnet1, CLRZ, PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP3 ( BFONET1, FNET4, CLK, CLRZ, PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP1 ( BFONET2, CLRZ, PREZ, BFONET1 ) ;


`endif

`ifdef TI_functiononly

	buf	TI_BUF_PRIM0 ( Q, BFONET1 ) ;

        buf #1 TI_BUF_PRIM1 ( QZ, BFONET2 ) ;


`else

           buf   TI_BUF_PRIM2 ( Q, BFONET1 ) ;
           buf   TI_BUF_PRIM3 ( QZ, BFONET2 ) ;
           not   TI_INV_PRIM3 ( QZ_NOT, QZ ) ; 
`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ , 1'b0 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND4 ( GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ , 1'b1 , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND5 ( GVC_Q_NOTEQ_DIN_CLRZ_NOT0_PREZ_NOT0_ , QZ_NOT , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND6 ( GVC_Q_NOT0_PREZ_NOT0_ , QZ_NOT , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND7 ( GVC_Q_NOT1_CLRZ_NOT0_ , QZ_NOT , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly


specify
    $recovery(posedge PREZ ,posedge CLRZ ,1 , GVCnotifier2_zd );
endspecify

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_DIN_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_;

    and TI_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_, GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_, GVC_Q_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_, GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_, GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ (TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_, GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_, GVC_Q_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_DIN_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_DIN_CLRZ_NOT0_PREZ_NOT0_, GVC_Q_NOTEQ_DIN_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ (TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_, GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_, TCHKON_NET);

`endif


specify
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ != 0  , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $setuphold(posedge PREZ &&& (TCHKON_NET != 0) , posedge CLRZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_PREZ_PREZ, GVC_CLRZ_CLRZ ); 
   $setuphold(posedge CLRZ &&& (TCHKON_NET != 0) , posedge PREZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_DIN_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_DIN_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ  &&& TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge PREZ  &&& TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

`endif // ifdef TETRAMAX
endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 09-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
// 12-jan-2010 Mazhar, Badarish: Updated to generate the new condition using
//             primary output (qz) for width check of clk (posedge and negedge)
//             Also for the above condition, D_OR_SD is replace by DIN.
// 13-jan-2010 Mazhar, Badarish: Reverted the changes done on 12-jan-2010, 
//             retaining only the update to use primary output QZ for width checks
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module SDB40 (CLK , CLRZ, D, PREZ, S, SD, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input PREZ;
   input S;
   input SD;
   output Q;
   output QZ;

`ifdef TETRAMAX
   _INV I1  ( CLRZ,CLR);
   _INV I2  ( PREZ,PRE);
   _NAND N1 ( CLR,PRE,CLR_PRE);
   _MUX M2  ( S, D, SD, DINT );
   _DFF FF1 ( !PREZ, !CLRZ, CLK, DINT, QINT);
   _INV I3  ( QINT,QZINT);
   _AND A1  ( CLRZ,QINT,Q1);
   _AND A2  ( PRE,CLR_PRE,Q2);
   _AND A3  ( QZINT,PREZ, Q3);
   _AND A4  ( CLR, CLR_PRE, Q4);
   _OR  O1  ( Q1,Q2,Q);
   _OR  O2  ( Q3,Q4,QZ);
`else
 


`ifdef TI_verilog    
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     parameter Xon = 1;
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_CLRZ_CLRZ  ,  GVC_PREZ_PREZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
        dlaudp   TI_DLA_UDP0 ( FNET4, DIN, IINVnet1, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP1 ( BFONET1, FNET4, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP0 ( BFONET2, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, BFONET1 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
        dlaudp   TI_DLA_UDP2 ( FNET4, DIN, IINVnet1, CLRZ, PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP3 ( BFONET1, FNET4, CLK, CLRZ, PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP1 ( BFONET2, CLRZ, PREZ, BFONET1 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          buf #1 TI_BUF_PRIM1 ( QZ, BFONET2 ) ;


`else

          buf  TI_BUF_PRIM2 ( Q, BFONET1 ) ;
          buf  TI_BUF_PRIM3 ( QZ, BFONET2 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ , 1'b0 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND4 ( GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ , 1'b1 , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND5 ( GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND6 ( GVC_Q_NOT0_PREZ_NOT0_ , Q , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND7 ( GVC_Q_NOT1_CLRZ_NOT0_ , Q , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly


specify
    $recovery(posedge PREZ ,posedge CLRZ ,1 , GVCnotifier2_zd );
endspecify

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_;

    and TI_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_, GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_, GVC_Q_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_, GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_, GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ (TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_, GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_, GVC_Q_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_, GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ (TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_, GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_, TCHKON_NET);

`endif


specify
      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ != 0  , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $setuphold(posedge PREZ &&& (TCHKON_NET != 0) , posedge CLRZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_PREZ_PREZ, GVC_CLRZ_CLRZ ); 
   $setuphold(posedge CLRZ &&& (TCHKON_NET != 0) , posedge PREZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ  &&& TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge PREZ  &&& TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

`endif // ifdef TETRAMAX
endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 09-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module SDB43 (CLK , CLRZ, D, PREZ, S, SD, Q ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input PREZ;
   input S;
   input SD;
   output Q;

`ifdef TETRAMAX
   _INV I1  ( CLRZ,CLR);
   _INV I2  ( PREZ,PRE);
   _NAND N1 ( CLR,PRE,CLR_PRE);
   _MUX M2  ( S, D, SD, DINT );
   _DFF FF1 ( !PREZ, !CLRZ, CLK, DINT, QINT);
   _INV I3  ( QINT,QZINT);
   _AND A1  ( CLRZ,QINT,Q1);
   _AND A2  ( PRE,CLR_PRE,Q2);
   _AND A3  ( QZINT,PREZ, Q3);
   _AND A4  ( CLR, CLR_PRE, Q4);
   _OR  O1  ( Q1,Q2,Q);
`else
 


`ifdef TI_verilog    
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     parameter Xon = 1;
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_CLRZ_CLRZ  ,  GVC_PREZ_PREZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
        dlaudp   TI_DLA_UDP0 ( FNET4, DIN, IINVnet1, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP1 ( BFONET1, FNET4, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP0 ( BFONET2, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, BFONET1 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
        dlaudp   TI_DLA_UDP2 ( FNET4, DIN, IINVnet1, CLRZ, PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP3 ( BFONET1, FNET4, CLK, CLRZ, PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP1 ( BFONET2, CLRZ, PREZ, BFONET1 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          buf  TI_BUF_PRIM1 ( QZ, BFONET2 ) ;


`else

          buf  TI_BUF_PRIM2 ( Q, BFONET1 ) ;
          buf  TI_BUF_PRIM3 ( QZ, BFONET2 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ , 1'b0 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND4 ( GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ , 1'b1 , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND5 ( GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND6 ( GVC_Q_NOT0_PREZ_NOT0_ , Q , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND7 ( GVC_Q_NOT1_CLRZ_NOT0_ , Q , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly


specify
    $recovery(posedge PREZ ,posedge CLRZ ,1 , GVCnotifier2_zd );
endspecify

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_;

    and TI_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_, GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_, GVC_Q_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_, GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_, GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ (TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_, GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_, GVC_Q_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_, GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ (TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_, GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_, TCHKON_NET);

`endif


specify
      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ != 0  , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $setuphold(posedge PREZ &&& (TCHKON_NET != 0) , posedge CLRZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_PREZ_PREZ, GVC_CLRZ_CLRZ ); 
   $setuphold(posedge CLRZ &&& (TCHKON_NET != 0) , posedge PREZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ  &&& TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge PREZ  &&& TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

`endif // ifdef TETRAMAX
endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 09-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module SDB44 (CLK , CLRZ, D, PREZ, S, SD,  QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input PREZ;
   input S;
   input SD;
   output QZ;

`ifdef TETRAMAX
   _INV I1  ( CLRZ,CLR);
   _INV I2  ( PREZ,PRE);
   _NAND N1 ( CLR,PRE,CLR_PRE);
   _MUX M2  ( S, D, SD, DINT );
   _DFF FF1 ( !PREZ, !CLRZ, CLK, DINT, QINT);
   _INV I3  ( QINT,QZINT);
   _AND A1  ( CLRZ,QINT,Q1);
   _AND A2  ( PRE,CLR_PRE,Q2);
   _AND A3  ( QZINT,PREZ, Q3);
   _AND A4  ( CLR, CLR_PRE, Q4);
   _OR  O2  ( Q3,Q4,QZ);
`else
 


`ifdef TI_verilog    
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     parameter Xon = 1;
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_CLRZ_CLRZ  ,  GVC_PREZ_PREZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
        dlaudp   TI_DLA_UDP0 ( FNET4, DIN, IINVnet1, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP1 ( BFONET1, FNET4, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP0 ( BFONET2, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ, BFONET1 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
        dlaudp   TI_DLA_UDP2 ( FNET4, DIN, IINVnet1, CLRZ, PREZ, GVCnotifier1 ) ;
        dlaudp   TI_DLA_UDP3 ( BFONET1, FNET4, CLK, CLRZ, PREZ, GVCnotifier2 ) ;
      dffqzudp   TI_QZ_UDP1 ( BFONET2, CLRZ, PREZ, BFONET1 ) ;


`endif

`ifdef TI_functiononly

	buf	TI_BUF_PRIM0 ( Q, BFONET1 ) ;

        buf #1 TI_BUF_PRIM1 ( QZ, BFONET2 ) ;


`else

           buf   TI_BUF_PRIM2 ( Q, BFONET1 ) ;
           buf   TI_BUF_PRIM3 ( QZ, BFONET2 ) ;
           not   TI_INV_PRIM3 ( QZ_NOT, QZ ) ; 
`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ , 1'b0 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND4 ( GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ , 1'b1 , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND5 ( GVC_Q_NOTEQ_DIN_CLRZ_NOT0_PREZ_NOT0_ , QZ_NOT , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND6 ( GVC_Q_NOT0_PREZ_NOT0_ , QZ_NOT , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND7 ( GVC_Q_NOT1_CLRZ_NOT0_ , QZ_NOT , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly


specify
    $recovery(posedge PREZ ,posedge CLRZ ,1 , GVCnotifier2_zd );
endspecify

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_DIN_CLRZ_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_;

    and TI_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_, GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_, GVC_Q_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_, GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_, GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ (TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_, GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_, GVC_Q_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_DIN_CLRZ_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_DIN_CLRZ_NOT0_PREZ_NOT0_, GVC_Q_NOTEQ_DIN_CLRZ_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ (TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_, GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_, TCHKON_NET);

`endif


specify
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_PREZ_NOT0_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_CLRZ_NOT0_ != 0  , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $setuphold(posedge PREZ &&& (TCHKON_NET != 0) , posedge CLRZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_PREZ_PREZ, GVC_CLRZ_CLRZ ); 
   $setuphold(posedge CLRZ &&& (TCHKON_NET != 0) , posedge PREZ,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier2_zd ,,, GVC_CLRZ_CLRZ, GVC_PREZ_PREZ ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_DIN_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_DIN_CLRZ_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ  &&& TCHKON_AND_GVC_Q_NOT0_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge PREZ  &&& TCHKON_AND_GVC_Q_NOT1_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

`endif // ifdef TETRAMAX
endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 09-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
// 12-jan-2010 Mazhar, Badarish: Updated to generate the new condition using
//             primary output (qz) for width check of clk (posedge and negedge)
//             Also for the above condition, D_OR_SD is replace by DIN.
// 13-jan-2010 Mazhar, Badarish: Reverted the changes done on 12-jan-2010, 
//             retaining only the update to use primary output QZ for width checks
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module SDC20 (CLK , CLRZ, D, S, SD, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input S;
   input SD;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_CLRZ_CLRZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, DIN, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, DIN, IINVnet1, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( BFONET1, FNET2, CLK, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_CLRZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_CLRZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_CLRZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT0_D_NOT0_S_WHATEVER_ , 1'b0 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;
    cons_udp TI_COND4 ( GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_;
    wire TCHKON_AND_Q;
    wire TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_;

    and TI_AND_GVC_S_NOT0_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_, GVC_S_NOT0_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ (TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_, GVC_SD_NOT0_D_NOT0_S_WHATEVER_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_, GVC_D_NOTEQ_SD_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_, GVC_S_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_, GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_, TCHKON_NET);

`endif


specify

      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& TCHKON_AND_Q != 0  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.3 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module SDC21 (CLK , CLRZ, D, LD, S, SD, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input LD;
   input S;
   input SD;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_CLRZ_CLRZ  ,  GVC_LD_LD  ; 

           not   TI_NOT_PRIM0 ( NOT_GVC_LD_LD, GVC_LD_LD ) ;
        mu1udp   TI_MUX2_UDP0 ( E2EG_6015, NOT_GVC_LD_LD, GVC_D_D, BFONET1 ) ;
        mu1udp   TI_MUX2_UDP1 ( DIN2, GVC_S_S, E2EG_6015, GVC_SD_SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, GVC_CLK_CLK ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, DIN2, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM2 ( NOT_LD, LD ) ;
        mu1udp   TI_MUX2_UDP2 ( E2EG_6015, NOT_LD, D, BFONET1 ) ;
        mu1udp   TI_MUX2_UDP3 ( DIN2, S, E2EG_6015, SD ) ;
           not   TI_NOT_PRIM3 ( IINVnet1, CLK ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, DIN2, IINVnet1, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( BFONET1, FNET2, CLK, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM4 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM5 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM6 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM7 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog
 
//  Logic enabling constraint check statements for verilog/verifault
 
  //  not TI_NOT_PRIM4 ( NOTENZ, GVC_ENZ_ENZ ) ;
    mu1udp   TI_MUX2_UDP4 ( DORQ_1, NOT_GVC_LD_LD, GVC_D_D, Q ) ;

    buf TI_BUF_PRIM3 ( DORQ , DORQ_1 ) ;
    not TI_NOT_PRIM5 ( NOTS, GVC_S_S ) ;
 
    and TI_AND_PRIM0 ( GVC_S_NOT1_LD_NOT0_CLRZ_NOT0_ , NOTS , GVC_LD_LD , GVC_CLRZ_CLRZ ) ;
    cons_udp TI_COND0 ( GVC_DORQ_NOTEQ_SD_CLRZ_NOT0_ , DORQ , GVC_SD_SD , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;
    and TI_AND_PRIM1 ( GVC_S_NOT0_CLRZ_NOT0_ , GVC_S_S , GVC_CLRZ_CLRZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_Q_S_NOT1_CLRZ_NOT0_ , Q, GVC_D_D, 1'b0, 1'b1, GVC_CLRZ_CLRZ , NOTS ) ;
    cons_udp TI_COND2 ( GVC_SD_NOT0_D_NOT0_S_WHATEVER_ , 1'b0 , GVC_SD_SD , DORQ , GVC_S_S , 1'b1 , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ , Q , GVC_SD_SD , DORQ , GVC_S_S , GVC_CLRZ_CLRZ , 1'b1 ) ;
 
`endif

`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_;
    wire TCHKON_AND_Q;
    wire TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_;
    wire TCHKON_AND_GVC_D_NOTEQ_Q_S_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_DORQ_NOTEQ_SD_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT1_LD_NOT0_CLRZ_NOT0_;

    and TI_AND_GVC_S_NOT0_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_, GVC_S_NOT0_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ (TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_, GVC_SD_NOT0_D_NOT0_S_WHATEVER_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_Q_S_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_Q_S_NOT1_CLRZ_NOT0_, GVC_D_NOTEQ_Q_S_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_, GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_DORQ_NOTEQ_SD_CLRZ_NOT0_ (TCHKON_AND_GVC_DORQ_NOTEQ_SD_CLRZ_NOT0_, GVC_DORQ_NOTEQ_SD_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT1_LD_NOT0_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_LD_NOT0_CLRZ_NOT0_, GVC_S_NOT1_LD_NOT0_CLRZ_NOT0_, TCHKON_NET);

`endif


specify

      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, ( TCHKON_AND_GVC_S_NOT1_LD_NOT0_CLRZ_NOT0_ != 0 ) , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, ( TCHKON_AND_GVC_S_NOT1_LD_NOT0_CLRZ_NOT0_ != 0 ) , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, ( TCHKON_AND_GVC_DORQ_NOTEQ_SD_CLRZ_NOT0_ != 0 ), GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, ( TCHKON_AND_GVC_DORQ_NOTEQ_SD_CLRZ_NOT0_ != 0 ), GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, ( TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0 ) , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, ( TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0 ) , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ != 0), GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $setuphold(posedge CLK,  posedge LD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, ( TCHKON_AND_GVC_D_NOTEQ_Q_S_NOT1_CLRZ_NOT0_ != 0 ), GVC_CLK_CLK, GVC_LD_LD ); 
   $setuphold(posedge CLK,  negedge LD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, ( TCHKON_AND_GVC_D_NOTEQ_Q_S_NOT1_CLRZ_NOT0_ != 0 ), GVC_CLK_CLK, GVC_LD_LD ); 
   $width(posedge CLK  &&& ( TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0 )  ,0.01 : 0.01 : 0.01 ,  0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& ( TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0 )  ,0.01 : 0.01 : 0.01 ,  0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& ( TCHKON_AND_Q != 0 )  ,0.01 : 0.01 : 0.01 ,  0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.3  05-Sep-2001 Removed the Copyright block
// v1.2  18-Sep-1999 Duplicate instance names were corrected
// v1.1  03-Sep-1999 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
// 13-jan-2010 Mazhar, Badarish: Updated to use primary output Q for
//             constraints check
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module SDC23 (CLK , CLRZ, D, S, SD, Q ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input S;
   input SD;
   output Q;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_CLRZ_CLRZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, DIN, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, DIN, IINVnet1, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( BFONET1, FNET2, CLK, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_CLRZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_CLRZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_CLRZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT0_D_NOT0_S_WHATEVER_ , 1'b0 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;
    cons_udp TI_COND4 ( GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_;
    wire TCHKON_AND_Q;
    wire TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_;

    and TI_AND_GVC_S_NOT0_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_, GVC_S_NOT0_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ (TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_, GVC_SD_NOT0_D_NOT0_S_WHATEVER_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_, GVC_D_NOTEQ_SD_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_, GVC_S_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_, GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_, TCHKON_NET);

`endif


specify

      (CLK  *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& TCHKON_AND_Q != 0  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module SDC24 (CLK , CLRZ, D, S, SD, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input S;
   input SD;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_CLRZ_CLRZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, DIN, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( Q, FNET2, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, DIN, IINVnet1, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( Q, FNET2, CLK, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          not #1 TI_NOT_PRIM2 ( QZ, Q ) ;


`else

          not  TI_NOT_PRIM3 ( QZ, Q ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_CLRZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_CLRZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_CLRZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT0_D_NOT0_S_WHATEVER_ , 1'b0 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;
    not TI_NOT_PRIM4 (GVCnet0 , GVC_SD_SD);
    not TI_NOT_PRIM5 (GVCnet1 , GVC_D_D);

   cons_udp TI_COND4 ( GVC_QZ_NOTEQ_SD_OR_D_CLRZ_NOT0_ , QZ , GVCnet0 , GVCnet1 , GVC_S_S , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_;

    and TI_AND_GVC_S_NOT0_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_, GVC_S_NOT0_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ (TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_, GVC_SD_NOT0_D_NOT0_S_WHATEVER_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_, GVC_D_NOTEQ_SD_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_QZ_NOTEQ_SD_OR_D_CLRZ_NOT0_ (TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_CLRZ_NOT0_, GVC_QZ_NOTEQ_SD_OR_D_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_, GVC_S_NOT1_CLRZ_NOT0_, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_QZ;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_QZ (NOT_TCHKON_OR_QZ, QZ, TCHKON_INV);

`endif


specify

      (CLK  *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& NOT_TCHKON_OR_QZ != 1  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models
//v2.0 12-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed

//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module SDC40 (CLK , CLRZ, D, S, SD, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input S;
   input SD;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_CLRZ_CLRZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, DIN, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, DIN, IINVnet1, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( BFONET1, FNET2, CLK, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_CLRZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_CLRZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_CLRZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT0_D_NOT0_S_WHATEVER_ , 1'b0 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;
    cons_udp TI_COND4 ( GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_;
    wire TCHKON_AND_Q;
    wire TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_;

    and TI_AND_GVC_S_NOT0_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_, GVC_S_NOT0_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ (TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_, GVC_SD_NOT0_D_NOT0_S_WHATEVER_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_, GVC_D_NOTEQ_SD_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_, GVC_S_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_, GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_, TCHKON_NET);

`endif


specify

      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& TCHKON_AND_Q != 0  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.3 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module SDC41 (CLK , CLRZ, D, LD, S, SD, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input LD;
   input S;
   input SD;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_CLRZ_CLRZ  ,  GVC_LD_LD  ; 

           not   TI_NOT_PRIM0 ( NOT_GVC_LD_LD, GVC_LD_LD ) ;
        mu1udp   TI_MUX2_UDP0 ( E2EG_6015, NOT_GVC_LD_LD, GVC_D_D, BFONET1 ) ;
        mu1udp   TI_MUX2_UDP1 ( DIN2, GVC_S_S, E2EG_6015, GVC_SD_SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, GVC_CLK_CLK ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, DIN2, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

           not   TI_NOT_PRIM2 ( NOT_LD, LD ) ;
        mu1udp   TI_MUX2_UDP2 ( E2EG_6015, NOT_LD, D, BFONET1 ) ;
        mu1udp   TI_MUX2_UDP3 ( DIN2, S, E2EG_6015, SD ) ;
           not   TI_NOT_PRIM3 ( IINVnet1, CLK ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, DIN2, IINVnet1, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( BFONET1, FNET2, CLK, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM4 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM5 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM6 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM7 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog
 
//  Logic enabling constraint check statements for verilog/verifault
 
  //  not TI_NOT_PRIM4 ( NOTENZ, GVC_ENZ_ENZ ) ;
    mu1udp   TI_MUX2_UDP4 ( DORQ_1, NOT_GVC_LD_LD, GVC_D_D, Q ) ;

    buf TI_BUF_PRIM3 ( DORQ , DORQ_1 ) ;
    not TI_NOT_PRIM5 ( NOTS, GVC_S_S ) ;
 
    and TI_AND_PRIM0 ( GVC_S_NOT1_LD_NOT0_CLRZ_NOT0_ , NOTS , GVC_LD_LD , GVC_CLRZ_CLRZ ) ;
    cons_udp TI_COND0 ( GVC_DORQ_NOTEQ_SD_CLRZ_NOT0_ , DORQ , GVC_SD_SD , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;
    and TI_AND_PRIM1 ( GVC_S_NOT0_CLRZ_NOT0_ , GVC_S_S , GVC_CLRZ_CLRZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_Q_S_NOT1_CLRZ_NOT0_ , Q, GVC_D_D, 1'b0, 1'b1, GVC_CLRZ_CLRZ , NOTS ) ;
    cons_udp TI_COND2 ( GVC_SD_NOT0_D_NOT0_S_WHATEVER_ , 1'b0 , GVC_SD_SD , DORQ , GVC_S_S , 1'b1 , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ , Q , GVC_SD_SD , DORQ , GVC_S_S , GVC_CLRZ_CLRZ , 1'b1 ) ;
 
`endif

`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_;
    wire TCHKON_AND_Q;
    wire TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_;
    wire TCHKON_AND_GVC_D_NOTEQ_Q_S_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_DORQ_NOTEQ_SD_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT1_LD_NOT0_CLRZ_NOT0_;

    and TI_AND_GVC_S_NOT0_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_, GVC_S_NOT0_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ (TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_, GVC_SD_NOT0_D_NOT0_S_WHATEVER_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_Q_S_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_Q_S_NOT1_CLRZ_NOT0_, GVC_D_NOTEQ_Q_S_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_, GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_DORQ_NOTEQ_SD_CLRZ_NOT0_ (TCHKON_AND_GVC_DORQ_NOTEQ_SD_CLRZ_NOT0_, GVC_DORQ_NOTEQ_SD_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT1_LD_NOT0_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_LD_NOT0_CLRZ_NOT0_, GVC_S_NOT1_LD_NOT0_CLRZ_NOT0_, TCHKON_NET);

`endif


specify

      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, ( TCHKON_AND_GVC_S_NOT1_LD_NOT0_CLRZ_NOT0_ != 0 ) , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, ( TCHKON_AND_GVC_S_NOT1_LD_NOT0_CLRZ_NOT0_ != 0 ) , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, ( TCHKON_AND_GVC_DORQ_NOTEQ_SD_CLRZ_NOT0_ != 0 ), GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, ( TCHKON_AND_GVC_DORQ_NOTEQ_SD_CLRZ_NOT0_ != 0 ), GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, ( TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0 ) , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, ( TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0 ) , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,( TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ != 0), GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $setuphold(posedge CLK,  posedge LD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, ( TCHKON_AND_GVC_D_NOTEQ_Q_S_NOT1_CLRZ_NOT0_ != 0 ), GVC_CLK_CLK, GVC_LD_LD ); 
   $setuphold(posedge CLK,  negedge LD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,, ( TCHKON_AND_GVC_D_NOTEQ_Q_S_NOT1_CLRZ_NOT0_ != 0 ), GVC_CLK_CLK, GVC_LD_LD ); 
   $width(posedge CLK  &&& ( TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0 )  ,0.01 : 0.01 : 0.01 ,  0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& ( TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0 )  ,0.01 : 0.01 : 0.01 ,  0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& ( TCHKON_AND_Q != 0 )  ,0.01 : 0.01 : 0.01 ,  0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.3  05-Sep-2001 Removed the Copyright block
// v1.2  18-Sep-1999 Duplicate instance names were corrected
// v1.1  03-Sep-1999 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
// 13-jan-2010 Mazhar, Badarish: Updated to use primary output Q for
//             constraints check
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module SDC43 (CLK , CLRZ, D, S, SD, Q ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input S;
   input SD;
   output Q;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_CLRZ_CLRZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, DIN, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, DIN, IINVnet1, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( BFONET1, FNET2, CLK, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_CLRZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_CLRZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_CLRZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT0_D_NOT0_S_WHATEVER_ , 1'b0 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;
    cons_udp TI_COND4 ( GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_;
    wire TCHKON_AND_Q;
    wire TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_;

    and TI_AND_GVC_S_NOT0_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_, GVC_S_NOT0_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ (TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_, GVC_SD_NOT0_D_NOT0_S_WHATEVER_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_, GVC_D_NOTEQ_SD_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_, GVC_S_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_, GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_, TCHKON_NET);

`endif


specify

      (CLK  *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& TCHKON_AND_Q != 0  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module SDC44 (CLK , CLRZ, D, S, SD, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input S;
   input SD;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_CLRZ_CLRZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, DIN, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( Q, FNET2, GVC_CLK_CLK, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, DIN, IINVnet1, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( Q, FNET2, CLK, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          not #1 TI_NOT_PRIM2 ( QZ, Q ) ;


`else

          not  TI_NOT_PRIM3 ( QZ, Q ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_CLRZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_CLRZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_CLRZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT0_D_NOT0_S_WHATEVER_ , 1'b0 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;
    not TI_NOT_PRIM4 (GVCnet0 , GVC_SD_SD);
    not TI_NOT_PRIM5 (GVCnet1 , GVC_D_D);

   cons_udp TI_COND4 ( GVC_QZ_NOTEQ_SD_OR_D_CLRZ_NOT0_ , QZ , GVCnet0 , GVCnet1 , GVC_S_S , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_;

    and TI_AND_GVC_S_NOT0_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_, GVC_S_NOT0_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ (TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_, GVC_SD_NOT0_D_NOT0_S_WHATEVER_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_, GVC_D_NOTEQ_SD_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_QZ_NOTEQ_SD_OR_D_CLRZ_NOT0_ (TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_CLRZ_NOT0_, GVC_QZ_NOTEQ_SD_OR_D_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_, GVC_S_NOT1_CLRZ_NOT0_, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_QZ;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_QZ (NOT_TCHKON_OR_QZ, QZ, TCHKON_INV);

`endif


specify

      (CLK  *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge CLRZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& NOT_TCHKON_OR_QZ != 1  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models
//v2.0 12-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed

//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module SDN20 (CLK , D, S, SD, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input S;
   input SD;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_nudp   TI_LACTHN_UDP0 ( FNET2, DIN, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_nudp   TI_LACTHN_UDP2 ( FNET2, DIN, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP3 ( BFONET1, FNET2, CLK, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_D_NOTEQ_SD_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , 1'b1 , 1'b1 ) ;
    cons_udp TI_COND1 ( GVC_Q_NOTEQ_SD_OR_D_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_D_NOTEQ_SD_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_;
    wire TCHKON_AND_S;
    wire TCHKON_AND_GVC_S_S;

    and TI_AND_GVC_D_NOTEQ_SD_ (TCHKON_AND_GVC_D_NOTEQ_SD_, GVC_D_NOTEQ_SD_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_, GVC_Q_NOTEQ_SD_OR_D_, TCHKON_NET);
    and TI_AND_S (TCHKON_AND_S, S, TCHKON_NET);
    and TI_AND_GVC_S_S (TCHKON_AND_GVC_S_S, GVC_S_S, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_S;
    wire NOT_TCHKON_OR_GVC_S_S;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_S (NOT_TCHKON_OR_S, S, TCHKON_INV);
    or TI_OR_GVC_S_S (NOT_TCHKON_OR_GVC_S_S, GVC_S_S, TCHKON_INV);

`endif


specify

      ( CLK *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      ( CLK *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_S_S != 1 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_S_S != 1 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_S != 0 , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_S != 0 , GVC_CLK_CLK, GVC_SD_SD ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.3 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module SDN21 (CLK , D, S, SD, Q ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input S;
   input SD;
   output Q;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_nudp   TI_LACTHN_UDP0 ( FNET2, DIN, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_nudp   TI_LACTHN_UDP2 ( FNET2, DIN, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP3 ( BFONET1, FNET2, CLK, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_D_NOTEQ_SD_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , 1'b1 , 1'b1 ) ;
    cons_udp TI_COND1 ( GVC_Q_NOTEQ_SD_OR_D_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_D_NOTEQ_SD_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_;
    wire TCHKON_AND_S;
    wire TCHKON_AND_GVC_S_S;

    and TI_AND_GVC_D_NOTEQ_SD_ (TCHKON_AND_GVC_D_NOTEQ_SD_, GVC_D_NOTEQ_SD_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_, GVC_Q_NOTEQ_SD_OR_D_, TCHKON_NET);
    and TI_AND_S (TCHKON_AND_S, S, TCHKON_NET);
    and TI_AND_GVC_S_S (TCHKON_AND_GVC_S_S, GVC_S_S, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_S;
    wire NOT_TCHKON_OR_GVC_S_S;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_S (NOT_TCHKON_OR_S, S, TCHKON_INV);
    or TI_OR_GVC_S_S (NOT_TCHKON_OR_GVC_S_S, GVC_S_S, TCHKON_INV);

`endif


specify

      (CLK *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_S_S != 1 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_S_S != 1 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_S != 0 , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_S != 0 , GVC_CLK_CLK, GVC_SD_SD ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.

// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version


//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module SDN22 (CLK , D, S, SD, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input S;
   input SD;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_nudp   TI_LACTHN_UDP0 ( FNET2, DIN, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP1 ( Q, FNET2, GVC_CLK_CLK, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_nudp   TI_LACTHN_UDP2 ( FNET2, DIN, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP3 ( Q, FNET2, CLK, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          not #1 TI_NOT_PRIM2 ( QZ, Q ) ;


`else

          not  TI_NOT_PRIM3 ( QZ, Q ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_D_NOTEQ_SD_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , 1'b1 , 1'b1 ) ;
    not TI_NOT_PRIM4 (GVCnet0 , GVC_SD_SD);
    not TI_NOT_PRIM5 (GVCnet1 , GVC_D_D);
    cons_udp TI_COND1 ( GVC_QZ_NOTEQ_SD_OR_D_ , QZ , GVCnet0 , GVCnet1 , GVC_S_S , 1'b1 , 1'b1 ) ;

`endif


`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_D_NOTEQ_SD_;
    wire TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_;
    wire TCHKON_AND_S;
    wire TCHKON_AND_GVC_S_S;

    and TI_AND_GVC_D_NOTEQ_SD_ (TCHKON_AND_GVC_D_NOTEQ_SD_, GVC_D_NOTEQ_SD_, TCHKON_NET);
    and TI_AND_GVC_QZ_NOTEQ_SD_OR_D_ (TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_, GVC_QZ_NOTEQ_SD_OR_D_, TCHKON_NET);
    and TI_AND_S (TCHKON_AND_S, S, TCHKON_NET);
    and TI_AND_GVC_S_S (TCHKON_AND_GVC_S_S, GVC_S_S, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_S;
    wire NOT_TCHKON_OR_GVC_S_S;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_S (NOT_TCHKON_OR_S, S, TCHKON_INV);
    or TI_OR_GVC_S_S (NOT_TCHKON_OR_GVC_S_S, GVC_S_S, TCHKON_INV);

`endif


specify

      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_S_S != 1 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_S_S != 1 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_S != 0 , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_S != 0 , GVC_CLK_CLK, GVC_SD_SD ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 09-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module SDN40 (CLK , D, S, SD, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input S;
   input SD;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_nudp   TI_LACTHN_UDP0 ( FNET2, DIN, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_nudp   TI_LACTHN_UDP2 ( FNET2, DIN, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP3 ( BFONET1, FNET2, CLK, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_D_NOTEQ_SD_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , 1'b1 , 1'b1 ) ;
    cons_udp TI_COND1 ( GVC_Q_NOTEQ_SD_OR_D_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_D_NOTEQ_SD_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_;
    wire TCHKON_AND_S;
    wire TCHKON_AND_GVC_S_S;

    and TI_AND_GVC_D_NOTEQ_SD_ (TCHKON_AND_GVC_D_NOTEQ_SD_, GVC_D_NOTEQ_SD_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_, GVC_Q_NOTEQ_SD_OR_D_, TCHKON_NET);
    and TI_AND_S (TCHKON_AND_S, S, TCHKON_NET);
    and TI_AND_GVC_S_S (TCHKON_AND_GVC_S_S, GVC_S_S, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_S;
    wire NOT_TCHKON_OR_GVC_S_S;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_S (NOT_TCHKON_OR_S, S, TCHKON_INV);
    or TI_OR_GVC_S_S (NOT_TCHKON_OR_GVC_S_S, GVC_S_S, TCHKON_INV);

`endif


specify

      ( CLK *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      ( CLK *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_S_S != 1 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_S_S != 1 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_S != 0 , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_S != 0 , GVC_CLK_CLK, GVC_SD_SD ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.3 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module SDN41 (CLK , D, S, SD, Q ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input S;
   input SD;
   output Q;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_nudp   TI_LACTHN_UDP0 ( FNET2, DIN, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_nudp   TI_LACTHN_UDP2 ( FNET2, DIN, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP3 ( BFONET1, FNET2, CLK, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_D_NOTEQ_SD_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , 1'b1 , 1'b1 ) ;
    cons_udp TI_COND1 ( GVC_Q_NOTEQ_SD_OR_D_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_D_NOTEQ_SD_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_;
    wire TCHKON_AND_S;
    wire TCHKON_AND_GVC_S_S;

    and TI_AND_GVC_D_NOTEQ_SD_ (TCHKON_AND_GVC_D_NOTEQ_SD_, GVC_D_NOTEQ_SD_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_, GVC_Q_NOTEQ_SD_OR_D_, TCHKON_NET);
    and TI_AND_S (TCHKON_AND_S, S, TCHKON_NET);
    and TI_AND_GVC_S_S (TCHKON_AND_GVC_S_S, GVC_S_S, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_S;
    wire NOT_TCHKON_OR_GVC_S_S;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_S (NOT_TCHKON_OR_S, S, TCHKON_INV);
    or TI_OR_GVC_S_S (NOT_TCHKON_OR_GVC_S_S, GVC_S_S, TCHKON_INV);

`endif


specify

      (CLK *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_S_S != 1 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_S_S != 1 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_S != 0 , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_S != 0 , GVC_CLK_CLK, GVC_SD_SD ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.

// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version


//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module SDN42 (CLK , D, S, SD, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input S;
   input SD;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_nudp   TI_LACTHN_UDP0 ( FNET2, DIN, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP1 ( Q, FNET2, GVC_CLK_CLK, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_nudp   TI_LACTHN_UDP2 ( FNET2, DIN, IINVnet1, GVCnotifier1 ) ;
       la_nudp   TI_LACTHN_UDP3 ( Q, FNET2, CLK, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          not #1 TI_NOT_PRIM2 ( QZ, Q ) ;


`else

          not  TI_NOT_PRIM3 ( QZ, Q ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_D_NOTEQ_SD_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , 1'b1 , 1'b1 ) ;
    not TI_NOT_PRIM4 (GVCnet0 , GVC_SD_SD);
    not TI_NOT_PRIM5 (GVCnet1 , GVC_D_D);
    cons_udp TI_COND1 ( GVC_QZ_NOTEQ_SD_OR_D_ , QZ , GVCnet0 , GVCnet1 , GVC_S_S , 1'b1 , 1'b1 ) ;

`endif


`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_D_NOTEQ_SD_;
    wire TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_;
    wire TCHKON_AND_S;
    wire TCHKON_AND_GVC_S_S;

    and TI_AND_GVC_D_NOTEQ_SD_ (TCHKON_AND_GVC_D_NOTEQ_SD_, GVC_D_NOTEQ_SD_, TCHKON_NET);
    and TI_AND_GVC_QZ_NOTEQ_SD_OR_D_ (TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_, GVC_QZ_NOTEQ_SD_OR_D_, TCHKON_NET);
    and TI_AND_S (TCHKON_AND_S, S, TCHKON_NET);
    and TI_AND_GVC_S_S (TCHKON_AND_GVC_S_S, GVC_S_S, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_S;
    wire NOT_TCHKON_OR_GVC_S_S;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_S (NOT_TCHKON_OR_S, S, TCHKON_INV);
    or TI_OR_GVC_S_S (NOT_TCHKON_OR_GVC_S_S, GVC_S_S, TCHKON_INV);

`endif


specify

      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_S_S != 1 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,NOT_TCHKON_OR_GVC_S_S != 1 , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_S != 0 , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_S != 0 , GVC_CLK_CLK, GVC_SD_SD ); 
   $width(posedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 09-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module SDP20 (CLK , D, PREZ, S, SD, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input PREZ;
   input S;
   input SD;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_PREZ_PREZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_pudp   TI_LACTHP_UDP0 ( FNET2, DIN, IINVnet1, GVC_PREZ_PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_PREZ_PREZ, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_pudp   TI_LACTHP_UDP2 ( FNET2, DIN, IINVnet1, PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP3 ( BFONET1, FNET2, CLK, PREZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_PREZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_PREZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT1_D_NOT1_S_WHATEVER_ , 1'b1 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;
    cons_udp TI_COND4 ( GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , GVC_PREZ_PREZ ) ;

`endif


`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_;
    wire TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_;

    and TI_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_ (TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_, GVC_SD_NOT1_D_NOT1_S_WHATEVER_, TCHKON_NET);
    and TI_AND_GVC_S_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_, GVC_S_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_, GVC_D_NOTEQ_SD_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_, GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT1_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_, GVC_S_NOT1_PREZ_NOT0_, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_Q;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_Q (NOT_TCHKON_OR_Q, Q, TCHKON_INV);

`endif


specify

      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_ != 0  , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge PREZ &&& NOT_TCHKON_OR_Q != 1  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.3 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module SDP23 (CLK , D, PREZ, S, SD, Q ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input PREZ;
   input S;
   input SD;
   output Q;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_PREZ_PREZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_pudp   TI_LACTHP_UDP0 ( FNET2, DIN, IINVnet1, GVC_PREZ_PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_PREZ_PREZ, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_pudp   TI_LACTHP_UDP2 ( FNET2, DIN, IINVnet1, PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP3 ( BFONET1, FNET2, CLK, PREZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;



`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_PREZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_PREZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT1_D_NOT1_S_WHATEVER_ , 1'b1 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;
    cons_udp TI_COND4 ( GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , GVC_PREZ_PREZ ) ;

`endif


`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_;
    wire TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_;

    and TI_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_ (TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_, GVC_SD_NOT1_D_NOT1_S_WHATEVER_, TCHKON_NET);
    and TI_AND_GVC_S_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_, GVC_S_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_, GVC_D_NOTEQ_SD_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_, GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT1_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_, GVC_S_NOT1_PREZ_NOT0_, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_Q;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_Q (NOT_TCHKON_OR_Q, Q, TCHKON_INV);

`endif


specify

      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_ != 0  , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge PREZ &&& NOT_TCHKON_OR_Q != 1  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 09-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module SDP24 (CLK , D, PREZ, S, SD, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input PREZ;
   input S;
   input SD;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_PREZ_PREZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_pudp   TI_LACTHP_UDP0 ( FNET2, DIN, IINVnet1, GVC_PREZ_PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_PREZ_PREZ, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_pudp   TI_LACTHP_UDP2 ( FNET2, DIN, IINVnet1, PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP3 ( BFONET1, FNET2, CLK, PREZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

	   buf	 TI_BUF_PRIM0 ( Q, BFONET1 ) ;

           not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

           buf   TI_BUF_PRIM1 ( Q, BFONET1 ) ;
           not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_PREZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_PREZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT1_D_NOT1_S_WHATEVER_ , 1'b1 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;
    not TI_NOT_PRIM4 (GVCnet0 , GVC_SD_SD);
    not TI_NOT_PRIM5 (GVCnet1 , GVC_D_D);
    cons_udp TI_COND4 ( GVC_QZ_NOTEQ_SD_OR_D_PREZ_NOT0_ , QZ , GVCnet0 , GVCnet1 , GVC_S_S , 1'b1 , GVC_PREZ_PREZ  ) ;

`endif


`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_;
    wire TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_;
    wire TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_PREZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_;

    and TI_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_ (TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_, GVC_SD_NOT1_D_NOT1_S_WHATEVER_, TCHKON_NET);
    and TI_AND_GVC_S_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_, GVC_S_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_, GVC_D_NOTEQ_SD_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_QZ_NOTEQ_SD_OR_D_PREZ_NOT0_ (TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_PREZ_NOT0_, GVC_QZ_NOTEQ_SD_OR_D_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT1_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_, GVC_S_NOT1_PREZ_NOT0_, TCHKON_NET);

   // wire TCHKON_INV;
    wire NOT_TCHKON_AND_Q;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

   // assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    and TI_AND_QZ (NOT_TCHKON_AND_QZ, QZ, TCHKON_NET);

`endif


specify

      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_ != 0  , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge PREZ &&& NOT_TCHKON_AND_QZ != 0  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.3 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module SDP40 (CLK , D, PREZ, S, SD, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input PREZ;
   input S;
   input SD;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_PREZ_PREZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_pudp   TI_LACTHP_UDP0 ( FNET2, DIN, IINVnet1, GVC_PREZ_PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_PREZ_PREZ, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_pudp   TI_LACTHP_UDP2 ( FNET2, DIN, IINVnet1, PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP3 ( BFONET1, FNET2, CLK, PREZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_PREZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_PREZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT1_D_NOT1_S_WHATEVER_ , 1'b1 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;
    cons_udp TI_COND4 ( GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , GVC_PREZ_PREZ ) ;

`endif


`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_;
    wire TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_;

    and TI_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_ (TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_, GVC_SD_NOT1_D_NOT1_S_WHATEVER_, TCHKON_NET);
    and TI_AND_GVC_S_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_, GVC_S_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_, GVC_D_NOTEQ_SD_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_, GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT1_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_, GVC_S_NOT1_PREZ_NOT0_, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_Q;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_Q (NOT_TCHKON_OR_Q, Q, TCHKON_INV);

`endif


specify

      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_ != 0  , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge PREZ &&& NOT_TCHKON_OR_Q != 1  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.3 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module SDP43 (CLK , D, PREZ, S, SD, Q ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input PREZ;
   input S;
   input SD;
   output Q;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_PREZ_PREZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_pudp   TI_LACTHP_UDP0 ( FNET2, DIN, IINVnet1, GVC_PREZ_PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_PREZ_PREZ, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_pudp   TI_LACTHP_UDP2 ( FNET2, DIN, IINVnet1, PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP3 ( BFONET1, FNET2, CLK, PREZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;



`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_PREZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_PREZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT1_D_NOT1_S_WHATEVER_ , 1'b1 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;
    cons_udp TI_COND4 ( GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , GVC_PREZ_PREZ ) ;

`endif


`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_;
    wire TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_;

    and TI_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_ (TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_, GVC_SD_NOT1_D_NOT1_S_WHATEVER_, TCHKON_NET);
    and TI_AND_GVC_S_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_, GVC_S_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_, GVC_D_NOTEQ_SD_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_, GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT1_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_, GVC_S_NOT1_PREZ_NOT0_, TCHKON_NET);

    wire TCHKON_INV;
    wire NOT_TCHKON_OR_Q;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

    assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    or TI_OR_Q (NOT_TCHKON_OR_Q, Q, TCHKON_INV);

`endif


specify

      (CLK *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> Q ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_ != 0  , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge PREZ &&& NOT_TCHKON_OR_Q != 1  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif


// Revision history:
// ----------------

//v1.1 09-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


 

module SDP44 (CLK , D, PREZ, S, SD, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input D;
   input PREZ;
   input S;
   input SD;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect
     wire GVCnotifier1;
     wire GVCnotifier2;


//  Verilog Notifier declaration section

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_PREZ_PREZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
       la_pudp   TI_LACTHP_UDP0 ( FNET2, DIN, IINVnet1, GVC_PREZ_PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP1 ( BFONET1, FNET2, GVC_CLK_CLK, GVC_PREZ_PREZ, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM1 ( IINVnet1, CLK ) ;
       la_pudp   TI_LACTHP_UDP2 ( FNET2, DIN, IINVnet1, PREZ, GVCnotifier1 ) ;
       la_pudp   TI_LACTHP_UDP3 ( BFONET1, FNET2, CLK, PREZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

	   buf	 TI_BUF_PRIM0 ( Q, BFONET1 ) ;

           not #1 TI_NOT_PRIM2 ( QZ, BFONET1 ) ;


`else

           buf   TI_BUF_PRIM1 ( Q, BFONET1 ) ;
           not  TI_NOT_PRIM3 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_PREZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_PREZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_PREZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , 1'b1 , GVC_PREZ_PREZ ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT1_D_NOT1_S_WHATEVER_ , 1'b1 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;
    not TI_NOT_PRIM4 (GVCnet0 , GVC_SD_SD);
    not TI_NOT_PRIM5 (GVCnet1 , GVC_D_D);
    cons_udp TI_COND4 ( GVC_QZ_NOTEQ_SD_OR_D_PREZ_NOT0_ , QZ , GVCnet0 , GVCnet1 , GVC_S_S , 1'b1 , GVC_PREZ_PREZ  ) ;

`endif


`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_;
    wire TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_;
    wire TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_PREZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_;

    and TI_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_ (TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_, GVC_SD_NOT1_D_NOT1_S_WHATEVER_, TCHKON_NET);
    and TI_AND_GVC_S_NOT0_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_, GVC_S_NOT0_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_, GVC_D_NOTEQ_SD_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_QZ_NOTEQ_SD_OR_D_PREZ_NOT0_ (TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_PREZ_NOT0_, GVC_QZ_NOTEQ_SD_OR_D_PREZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT1_PREZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_, GVC_S_NOT1_PREZ_NOT0_, TCHKON_NET);

   // wire TCHKON_INV;
    wire NOT_TCHKON_AND_Q;

    //not TI_NOT_TCHKON (TCHKON_INV, TCHKON);

   // assign TCHKON_INV = TCHKON ? 1'b0 : 1'b1 ;
    and TI_AND_QZ (NOT_TCHKON_AND_QZ, QZ, TCHKON_NET);

`endif


specify

      (CLK *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (PREZ *> QZ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);


`ifdef TI_verilog 

   $setuphold(posedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(posedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(posedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(posedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_PREZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge PREZ,  posedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT1_D_NOT1_S_WHATEVER_ != 0  , GVC_PREZ_PREZ , GVC_CLK_CLK);
   $width(posedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(negedge CLK  &&& TCHKON_AND_GVC_QZ_NOTEQ_SD_OR_D_PREZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge PREZ &&& NOT_TCHKON_AND_QZ != 0  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.3 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models

//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module SNC20 (CLK , CLRZ, D, S, SD, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input S;
   input SD;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect


//  Verilog Notifier declaration section

    wire GVCnotifier1 ;
    wire GVCnotifier2 ;

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_CLRZ_CLRZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
           not   TI_NOT_PRIM1 ( IINVnet2, IINVnet1 ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, DIN, IINVnet2, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, FNET2, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM2 ( IINVnet1, CLK ) ;
           not   TI_NOT_PRIM3 ( IINVnet2, IINVnet1 ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, DIN, IINVnet2, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( BFONET1, FNET2, IINVnet1, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM4 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM5 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_CLRZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_CLRZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_CLRZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT0_D_NOT0_S_WHATEVER_ , 1'b0 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;
    cons_udp TI_COND4 ( GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_;
    wire TCHKON_AND_Q;
    wire TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_;

    and TI_AND_GVC_S_NOT0_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_, GVC_S_NOT0_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ (TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_, GVC_SD_NOT0_D_NOT0_S_WHATEVER_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_, GVC_D_NOTEQ_SD_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_, GVC_S_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_, GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_, TCHKON_NET);

`endif


specify

      (CLK  *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK  *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(negedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(negedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(negedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(negedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(negedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(negedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge CLRZ,  negedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& TCHKON_AND_Q != 0  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

// 24 Apr 2006 : Sharavathi : Removed TI_veritime options and updated to support 
//                                Simulation without transimiting X when violation
//                                occurs by using Xon

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine



`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

// Verilog Interface section

module SNC40 (CLK , CLRZ, D, S, SD, Q, QZ ) ;

// Verilog Port Declaration section

   input CLK;
   input CLRZ;
   input D;
   input S;
   input SD;
   output Q;
   output QZ;


`ifdef TI_verilog    
    parameter Xon = 1;
    parameter TCHKON = 1;
    wire TCHKON_NET;
    assign TCHKON_NET = TCHKON ? 1'b1 : 1'b0 ;
//    buf TI_BUF_TCHKON (TCHKON_NET, TCHKON);
`endif

`ifdef TI_openhdl
`else
  `protect


//  Verilog Notifier declaration section

    wire GVCnotifier1 ;
    wire GVCnotifier2 ;

    reg GVCnotifier1_zd ;
    reg GVCnotifier2_zd ;

// Xon controlability

`ifdef TI_verilog
   and TI_GVCnotifier1 (GVCnotifier1, Xon, GVCnotifier1_zd);
   and TI_GVCnotifier2 (GVCnotifier2, Xon, GVCnotifier2_zd);
`endif 

// Verilog Structure section (in terms of gate prims)

 
`ifdef TI_verilog

// Net Declared for negative timing check
     wire  GVC_CLK_CLK ,  GVC_D_D  ,  GVC_S_S  ,  GVC_SD_SD  ,  GVC_CLRZ_CLRZ  ; 

        mu1udp   TI_MUX2_UDP0 ( DIN, GVC_S_S, GVC_D_D, GVC_SD_SD ) ;
           not   TI_NOT_PRIM0 ( IINVnet1, GVC_CLK_CLK ) ;
           not   TI_NOT_PRIM1 ( IINVnet2, IINVnet1 ) ;
       la_cudp   TI_LACTHC_UDP0 ( FNET2, DIN, IINVnet2, GVC_CLRZ_CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP1 ( BFONET1, FNET2, IINVnet1, GVC_CLRZ_CLRZ, GVCnotifier2 ) ;


`else

        mu1udp   TI_MUX2_UDP1 ( DIN, S, D, SD ) ;
           not   TI_NOT_PRIM2 ( IINVnet1, CLK ) ;
           not   TI_NOT_PRIM3 ( IINVnet2, IINVnet1 ) ;
       la_cudp   TI_LACTHC_UDP2 ( FNET2, DIN, IINVnet2, CLRZ, GVCnotifier1 ) ;
       la_cudp   TI_LACTHC_UDP3 ( BFONET1, FNET2, IINVnet1, CLRZ, GVCnotifier2 ) ;


`endif

`ifdef TI_functiononly

          buf #1 TI_BUF_PRIM0 ( Q, BFONET1 ) ;
          not #1 TI_NOT_PRIM4 ( QZ, BFONET1 ) ;


`else

          buf  TI_BUF_PRIM1 ( Q, BFONET1 ) ;
          not  TI_NOT_PRIM5 ( QZ, BFONET1 ) ;

`endif

`ifdef TI_verilog

//  Logic enabling constraint check statements for verilog/verifault

    cons_udp TI_COND0 ( GVC_S_NOT1_CLRZ_NOT0_ , GVC_S_S , 1'b1 , 1'b1 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND1 ( GVC_D_NOTEQ_SD_CLRZ_NOT0_ , GVC_D_D , GVC_SD_SD , 1'b0 , 1'b1 , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND2 ( GVC_S_NOT0_CLRZ_NOT0_ , GVC_S_S , 1'b0 , 1'b0 , 1'bx , GVC_CLRZ_CLRZ , 1'b1 ) ;
    cons_udp TI_COND3 ( GVC_SD_NOT0_D_NOT0_S_WHATEVER_ , 1'b0 , GVC_SD_SD , GVC_D_D , GVC_S_S , 1'b1 , 1'b1 ) ;
    cons_udp TI_COND4 ( GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ , Q , GVC_SD_SD , GVC_D_D , GVC_S_S , GVC_CLRZ_CLRZ , 1'b1 ) ;

`endif



`ifdef TI_functiononly

`else

`ifdef TI_verilog

    wire TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_;
    wire TCHKON_AND_Q;
    wire TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_;
    wire TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_;
    wire TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_;

    and TI_AND_GVC_S_NOT0_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_, GVC_S_NOT0_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_Q (TCHKON_AND_Q, Q, TCHKON_NET);
    and TI_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ (TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_, GVC_SD_NOT0_D_NOT0_S_WHATEVER_, TCHKON_NET);
    and TI_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ (TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_, GVC_D_NOTEQ_SD_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_S_NOT1_CLRZ_NOT0_ (TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_, GVC_S_NOT1_CLRZ_NOT0_, TCHKON_NET);
    and TI_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ (TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_, GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_, TCHKON_NET);

`endif


specify

      (CLK  *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLK  *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> Q  ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);
      (CLRZ *> QZ ) = (0.100000:0.100000:0.100000 , 0.100000:0.100000:0.100000);

`ifdef TI_verilog 

   $setuphold(negedge CLK,  posedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(negedge CLK,  negedge D,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT1_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_D_D ); 
   $setuphold(negedge CLK,  posedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(negedge CLK,  negedge S,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_D_NOTEQ_SD_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_S_S ); 
   $setuphold(negedge CLK,  posedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $setuphold(negedge CLK,  negedge SD,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_S_NOT0_CLRZ_NOT0_ != 0  , GVC_CLK_CLK, GVC_SD_SD ); 
   $recrem(posedge CLRZ,  negedge CLK,  0.01: 0.01: 0.01,  0.01: 0.01: 0.01, GVCnotifier1_zd ,,TCHKON_AND_GVC_SD_NOT0_D_NOT0_S_WHATEVER_ != 0  , GVC_CLRZ_CLRZ , GVC_CLK_CLK);
   $width(negedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 
   $width(posedge CLK  &&& TCHKON_AND_GVC_Q_NOTEQ_SD_OR_D_CLRZ_NOT0_ != 0   ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier1_zd) ; 
   $width(negedge CLRZ &&& TCHKON_AND_Q != 0  ,0.01 : 0.01 : 0.01 , 0 , GVCnotifier2_zd) ; 

`endif

endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------
// v1.4 08-Aug-2007 :Dundappa.
//                  Added the default delay of 1 for the output pins.
// v1.3  14-Jan-2002 Conditional paths have been modified in the specify section to
//                   take care of proper timing annotation Track Id 23313
// v1.2  05-Sep-2001 Removed the Copyright block
// v1.1  13-Dec-1998 Initial Version

// 24 Apr 2006 : Sharavathi : Removed TI_veritime options and updated to support 
//                                Simulation without transimiting X when violation
//                                occurs by using Xon

//v2.0 6-oct-2009 Mathangi Updated for non aligned models
//v2.0 9-Oct-2009 Mathangi removed "TI_veritime" defination from models
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module SPAREPOLYCAP11 () ;

endmodule
`endcelldefine







// Revision history:
// ----------------

//v1.0 16-May-2008 :Santosh: First version.
//v2.0 13-Oct-2009 :Mathangi: Updated delay mode distributed to 1ps/1ps from 1ns/1ns

//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module SPAREPOLYCAP16 () ;

endmodule
`endcelldefine







// Revision history:
// ----------------

//v1.0 16-May-2008 :Santosh: First version.
//v2.0 13-Oct-2009 :Mathangi: Updated delay mode distributed to 1ps/1ps from 1ns/1ns

//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module SPAREPOLYCAP32 () ;

endmodule
`endcelldefine







// Revision history:
// ----------------

//v1.0 16-May-2008 :Santosh: First version.
//v2.0 13-Oct-2009 :Mathangi: Updated delay mode distributed to 1ps/1ps from 1ns/1ns

//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module SPAREPOLYLDCAP11 () ;

endmodule
`endcelldefine







// Revision history:
// ----------------

//v1.0 16-May-2008 :Santosh: First version.
//v2.0 13-Oct-2009 :Mathangi: Updated delay mode distributed to 1ps/1ps from 1ns/1ns

//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module SPAREPOLYLDCAP16 () ;

endmodule
`endcelldefine







// Revision history:
// ----------------

//v1.0 16-May-2008 :Santosh: First version.
//v2.0 13-Oct-2009 :Mathangi: Updated delay mode distributed to 1ps/1ps from 1ns/1ns

//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine

`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module SPAREPOLYLDCAP32 () ;

endmodule
`endcelldefine







// Revision history:
// ----------------

//v1.0 16-May-2008 :Santosh: First version.
//v2.0 13-Oct-2009 :Mathangi: Updated delay mode distributed to 1ps/1ps from 1ns/1ns

`resetall
`ifdef TI_functiononly
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

primitive srudp_21
`protect
(q, s, r, nt);

input s, r, nt;
output q;
reg q;

table
//	s   r  nt  : q :	q;
      (?1)  1  ?   : ? :	1;
        1 (?1) ?   : ? :	1;
      (?1)  0  ?   : ? :	1;
	1 (?0) ?   : ? :	1;
      (?1)  x  ?   : ? :	1;
	1 (?x) ?   : ? :	1; 
      (?0)  1  ?   : ? :	0;
        0 (?1) ?   : ? :	0;
      (?0)  0  ?   : ? :	-;
	0 (?0) ?   : ? :	-;
       x (?0)  ?   : 1 :	1;
      (?x)  0  ?   : 1 :	1; 
      (?0)  x  ?   : 0 :	0;
	0 (?x) ?   : 0 :	0; 
	?  ?   *   : ? :	x;

endtable
`endprotect
endprimitive 

// 19 Dec 2006 : Sharavathi : changed the timescale for functiononly option to 
//                            1ns/1ps
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
`resetall
`ifdef TI_functiononly
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

primitive srudp
`protect
(q, s, r, nt);

input s, r, nt;
output q;
reg q;

table
//	s   r  nt  : q :	q;
  (?0)  0  ?   : ? :	0;
	0 (?0) ?   : ? :	0;
  (?1)  0  ?   : ? :	0;
	1 (?0) ?   : ? :	0;
  (?x)  0  ?   : ? :	0;
    x (?0) ?   : ? :	0;
  (?0)  1  ?   : ? :	1;
	0 (?1) ?   : ? :	1;
  (?1)  1  ?   : ? :	-;
	1 (?1) ?   : ? :	-;
  (?1)  x  ?   : 0 :	0;
	1 (?x) ?   : 0 :	0; 
  (?x)  1  ?   : 1 :    1;
    x (?1) ?   : 1 :    1;
	?  ?   *   : ? :	x;

endtable
`endprotect
endprimitive 

// 19 Dec 2006 : Sharavathi : changed the timescale for functiononly option to 
//                            1ns/1ps
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
`resetall
`ifdef TI_functiononly
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

primitive srudpz_21
`protect
(q, s, r, nt);

input s, r, nt;
output q;
reg q;

table

//	s   r  nt   :q: q;
      (?0)  0   ?   :?: -;
	0 (?0)  ?   :?: -;
      (?1)  0   ?   :?: 0;
        1 (?0)  ?   :?: 0;
      (?0)  1   ?   :?: 1;
	0  (?1) ?   :?: 1;
        x  (?1) ?   :?: 1;
      (?x)  1   ?   :?: 1;
      (?1)  1   ?   :?: 1;
	1  (?1) ?   :?: 1;
      (?0)  x   ?   :1: 1;
	0  (?x) ?   :1: 1;
      (?x)  0   ?   :0: 0;
        x (?0)  ?   :0: 0;
	?   ?   *   :?: x;

endtable
`endprotect
endprimitive 

// 19 Dec 2006 : Sharavathi : changed the timescale for functiononly option to 
//                            1ns/1ps
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
`resetall
`ifdef TI_functiononly
    `timescale 1ps / 1ps
`else
    `timescale 1ns / 1ps
`endif

primitive srudpz
`protect
(q, s, r, nt);

input s, r, nt;
output q;
reg q;

table

//	s   r  nt   :q: q;
  (?0)  0   ?   :?: 0;
	0 (?0)  ?   :?: 0;
  (?1)  0   ?   :?: 1;
    1  (?0) ?   :?: 1;
  (?0)  1   ?   :?: 0;
	0  (?1) ?   :?: 0;
  (?0)  x   ?   :?: 0;
    0  (?x) ?   :?: 0;
  (?1)  1   ?   :?: -;
	1  (?1) ?   :?: -;
  (?1)  x   ?   :1: 1;
	1  (?x) ?   :1: 1;
  (?x)  1   ?   :0: 0;
    x (?1)  ?   :0: 0;
	?   ?   *   :?: x;

endtable
`endprotect
endprimitive 

// 19 Dec 2006 : Sharavathi : changed the timescale for functiononly option to 
//                            1ns/1ps
//v2.0 9-oct-2009 Mathangi Updated for timescale 1ps/1ps for delay_mode_distributed
//---------------------------------------------------------------------
// Copyright (c) 2010 TEXAS INSTRUMENTS, Inc.                         
// All rights reserved                                                 
//                                                                     
// This is an UNPUBLISHED work created in the year stated above.       
// TEXAS INSTRUMENTS owns all rights in and to the work and intends to 
// maintain it and protect it as unpublished copyright. In the event   
// of either inadvertant or deliberate publication, the above stated   
// date shall be treated as the year of first publication. In the event
// of such publication, Texas Instruments intends to enforce its rights
// in the work under the copyright laws as a published work.           
//                                                                     
// These commodities are under U.S. Government distribution license    
// control. As such, they are not be re-exported without prior approval
// from the U.S. Department of Commerce.                               
//                                                                     
//---------------------------------------------------------------------

// Revision history:
// ----------------

`resetall
`ifdef TI_verifault
`suppress_faults
`enable_portfaults
`endif

`celldefine





`ifdef TI_functiononly
    `delay_mode_distributed
    `timescale 1ps / 1ps
`else
    `delay_mode_path
    `timescale 1ns / 1ps
`endif

// Verilog Interface section


module TO020 ( ZERO, ONE ) ;

// Verilog Port Declaration section
    output ZERO;
    output ONE;

`ifdef TI_openhdl
`else
  `protect

// Verilog Structure section (in terms of gate prims)

           buf #0 TI_BUF_PRIM0 (ONE, 1'b1) ;
           buf #0 TI_BUF_PRIM1 (ZERO, 1'b0) ;

`ifdef TI_functiononly
`else

specify


endspecify
`endif

  `endprotect
`endif

endmodule

`endcelldefine

`ifdef TI_verifault
`nosuppress_faults
`disable_portfaults
`endif

// Revision history:
// ----------------

//v1.1 08-Aug-2007 :Dundappa.
//                  Added the default delay of 0 for the output pins.

//v1.0 17-Aug-2005 :Verilog Port Declaration section:
//                  Change in the Port order, in sync with module defination
//V2.0 12-Oct-2009 :Updated time scale to 1ps/1ps

